/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   riscv_i32_alu.cdl
 * @brief  ALU for i32 RISC-V implementation
 *
 * CDL implementation of RISC-V i32 ALU based on the RISC-V
 * specification v2.1.
 *
 */

/*a Includes
 */
include "cpu/riscv/riscv_pipeline_types.h"
include "cpu/riscv/riscv_internal_types.h"
include "cpu/riscv/riscv.h"

/*a Constants
 */
constant integer coproc_force_disable=0;
constant integer debug_force_disable=0;

/*a Module
 */
module riscv_i32_pipeline_control_flow( input  t_riscv_pipeline_state        pipeline_state,
                                        input  t_riscv_fetch_req             ifetch_req,
                                        input  t_riscv_pipeline_response     pipeline_response,
                                        output t_riscv_pipeline_control      pipeline_control,
                                        input t_riscv_i32_coproc_response    coproc_response,
                                        output  t_riscv_mem_access_req       dmem_access_req,
                                        output  t_riscv_csr_access           csr_access,
                                        output t_riscv_i32_coproc_response   pipeline_coproc_response,
                                        output t_riscv_i32_coproc_controls   coproc_controls,
                                        output t_riscv_csr_controls          csr_controls,
                                        output t_riscv_i32_trace             trace,
                                        input  t_riscv_config                riscv_config
    )
"""

"""
{
    comb t_riscv_i32_control_data  control_data;
    comb t_riscv_i32_control_flow  control_flow;
    control_flow_code : {
        control_flow.trap = {*=0};
        control_flow.branch_taken = 0;
        control_flow.jalr = 0;
        control_flow.next_pc = 0;
        control_flow.trap.pc = control_data.pc;
        control_flow.async_cancel = 0;
        control_flow.trap.to_mode = pipeline_state.interrupt_to_mode;
        part_switch (control_data.idecode.op) {
        case riscv_op_branch:   { control_flow.branch_taken = pipeline_response.exec.branch_condition_met; }
        case riscv_op_jal:      { control_flow.branch_taken=1; }
        case riscv_op_jalr:     { control_flow.branch_taken=1; control_flow.jalr=1; }
        case riscv_op_system:   {
            if (control_data.idecode.subop==riscv_subop_mret) {
                control_flow.trap.ret = 1;
                control_flow.trap.cause = riscv_trap_cause_ret_mret;
            }
            if (control_data.idecode.subop==riscv_subop_ecall) {
                control_flow.trap.valid = 1;
                control_flow.trap.cause = riscv_trap_cause_mecall;
            }
            if (control_data.idecode.subop==riscv_subop_ebreak) {
                control_flow.trap.valid = 1;
                control_flow.trap.ebreak_to_dbg = pipeline_state.ebreak_to_dbg;
                control_flow.trap.cause = riscv_trap_cause_breakpoint;
                control_flow.trap.value = control_data.pc;
            }
        }
        }
        if (!control_data.exec_committed) {
            control_flow.trap.valid = 0;
            control_flow.trap.ret = 0;
            control_flow.trap.ebreak_to_dbg = 0;
            control_flow.branch_taken = 0;
        }
        
        if (control_data.valid && control_data.idecode.illegal) { // exec_committed will be zero
            control_flow.trap.valid = 1;
            control_flow.trap.ret = 0;
            control_flow.trap.cause = riscv_trap_cause_illegal_instruction;
            control_flow.trap.value = control_data.instruction_data;
        }
        if (control_data.valid && control_data.idecode.illegal_pc) { // exec_committed will be zero
            control_flow.trap.valid = 1;
            control_flow.trap.ret = 0;
            control_flow.trap.cause = riscv_trap_cause_instruction_misaligned;
            control_flow.trap.value = control_data.pc;
        }
        if (pipeline_state.interrupt_req && !pipeline_response.exec.interrupt_block) {
            control_flow.async_cancel = 1;
            control_flow.trap.valid = 1;
            control_flow.trap.ret = 0;
            control_flow.trap.cause = riscv_trap_cause_interrupt;
            control_flow.trap.cause[4;0] = pipeline_state.interrupt_number;
            control_flow.trap.value = control_data.pc;
        }
    }
    code : {

        control_data = {*=0};
        control_data = { instruction_data = pipeline_response.exec.instruction.data,
                                   pc               = pipeline_response.exec.pc,
                                   interrupt_ack    = 1,
                                   valid            = pipeline_response.exec.valid,
                         exec_committed   = pipeline_response.exec.valid && !pipeline_response.exec.cannot_start,
                                   idecode          = pipeline_response.exec.idecode,
                                   first_cycle = pipeline_response.exec.first_cycle
        };
        if (!pipeline_response.exec.valid) {
            control_data.pc = pipeline_response.decode.valid ? pipeline_response.decode.pc : pipeline_state.fetch_pc;
        }

        pipeline_control.valid = pipeline_state.valid;
        pipeline_control.fetch_action = pipeline_state.fetch_action;
        pipeline_control.fetch_pc = pipeline_state.fetch_pc;
        pipeline_control.mode = pipeline_state.mode;
        pipeline_control.error = pipeline_state.error;
        pipeline_control.tag = pipeline_state.tag;
        pipeline_control.halt = pipeline_state.halt;
        pipeline_control.interrupt_req = pipeline_state.interrupt_req;
        pipeline_control.interrupt_number = pipeline_state.interrupt_number;
        pipeline_control.ebreak_to_dbg = pipeline_state.ebreak_to_dbg;
        pipeline_control.interrupt_to_mode = pipeline_state.interrupt_to_mode;
        pipeline_control.instruction_data = pipeline_state.instruction_data;
        pipeline_control.instruction_debug = pipeline_state.instruction_debug;

        pipeline_control.async_cancel       = control_flow.async_cancel;
        pipeline_control.pc_if_mispredicted = control_flow.jalr ? pipeline_response.exec.branch_target : pipeline_response.exec.pc_if_mispredicted;
        pipeline_control.branch_taken       = control_flow.branch_taken;
        pipeline_control.jalr               = control_flow.jalr && (pipeline_response.exec.idecode.rs1!=0);
        pipeline_control.trap               = control_flow.trap;

        pipeline_coproc_response = coproc_response;
        if (coproc_force_disable || riscv_config.coproc_disable) {
            pipeline_coproc_response = {*=0};
        }

        pipeline_control.exec_cannot_start    = pipeline_response.exec.cannot_start     || pipeline_coproc_response.cannot_start;
        pipeline_control.exec_cannot_complete = pipeline_response.exec.cannot_complete  || pipeline_coproc_response.cannot_complete;
        if (pipeline_response.exec.first_cycle && pipeline_response.exec.valid && pipeline_control.exec_cannot_start) {
            pipeline_control.exec_cannot_complete = 1;
        }
        pipeline_control.exec_committed       = pipeline_response.exec.valid && !pipeline_control.exec_cannot_complete;
        pipeline_control.decode_cannot_complete = pipeline_response.decode.valid && pipeline_response.exec.valid && pipeline_control.exec_cannot_complete;

        dmem_access_req = pipeline_response.exec.dmem_access_req;
        if (!pipeline_control.exec_committed) { dmem_access_req.valid = 0; }

        csr_access = pipeline_response.exec.csr_access;
        if (!pipeline_response.exec.valid || pipeline_response.exec.idecode.illegal) {
            csr_access.access = riscv_csr_access_none;
        }
        csr_access.access_cancelled =  pipeline_control.async_cancel;



        //pipeline_control.alu_flush_pipeline     = ifetch_req.flush_pipeline;
        pipeline_control.flush_decode     = ifetch_req.flush_pipeline;
        pipeline_control.flush_fetch     = 0;
        pipeline_control.flush_exec     = 0;

        if (pipeline_response.exec.valid && (pipeline_control.branch_taken != pipeline_response.exec.predicted_branch)) {
            pipeline_control.flush_fetch     = 1;
            pipeline_control.flush_decode    = 1;
        }
        if (pipeline_control.trap.valid) {
            pipeline_control.flush_fetch     = 1;
            pipeline_control.flush_decode     = 1;
        }
        if (pipeline_control.trap.ret) {
            pipeline_control.flush_fetch     = 1;
            pipeline_control.flush_decode     = 1;
        }
        if (pipeline_state.instruction_debug.valid) {
            pipeline_control.flush_fetch     = 0;
        }

    }

    /*b CSR controls */
    csr_controls : {
        /*b CSR controls - post trap detection */
        csr_controls = {*=0};
        csr_controls.retire       = pipeline_response.exec.valid && pipeline_control.exec_committed;
        csr_controls.trap         = pipeline_control.trap;
    }

    /*b Coprocessor interface */
    coprocessor_interface """
    Drive the coprocessor controls unless disabled; mirror the pipeline combs

    Probably only legal if there is a decode stage - or if the coprocessor knows there is not
    """: {
        coproc_controls.dec_idecode        = pipeline_response.decode.idecode;
        coproc_controls.dec_idecode_valid  = pipeline_response.decode.valid && !pipeline_state.interrupt_req;
        coproc_controls.dec_to_alu_blocked = pipeline_response.exec.cannot_complete || coproc_response.cannot_complete;
        coproc_controls.alu_rs1 = pipeline_response.exec.rs1;
        coproc_controls.alu_rs2 = pipeline_response.exec.rs2;
        coproc_controls.alu_flush_pipeline  = pipeline_control.flush_decode; // pipeline_fetch_data.dec_flush_pipeline;
        coproc_controls.alu_cannot_start    = pipeline_response.exec.cannot_start    || coproc_response.cannot_start;
        coproc_controls.alu_cannot_complete = pipeline_response.exec.cannot_complete || coproc_response.cannot_complete;
        if (coproc_force_disable || riscv_config.coproc_disable) {
            coproc_controls = {*=0};
        }
    }

    /*b Trace */
    trace """
    Map the pipeline output to the trace
    """: {
        trace = {*=0};
        trace.instr_valid    = pipeline_response.exec.valid && pipeline_control.exec_committed;
        trace.instr_pc       = pipeline_response.exec.pc;
        trace.mode           = pipeline_state.mode;
        trace.instruction    = pipeline_response.exec.instruction.data;
        trace.rfw_retire     = pipeline_response.rfw.valid;
        trace.rfw_data_valid = pipeline_response.rfw.rd_written;
        trace.rfw_rd         = pipeline_response.rfw.rd;
        trace.rfw_data       = pipeline_response.rfw.data;
        trace.branch_taken   = pipeline_control.branch_taken;
        trace.trap           = pipeline_control.trap.valid;
        trace.ret            = pipeline_control.trap.ret;
        trace.jalr           = pipeline_control.jalr;
        trace.branch_target  = ifetch_req.address;
        trace.bkpt_valid     = 0;
        trace.bkpt_reason    = 0;
    }
}
