/** @copyright (C) 2019,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   gbe_axi4s32.cdl
 * @brief  GbE MAC (supporting 10/100/1000) full duplex using AXI-4S to GMII
 *
 * CDL implementation of a fully synchronous GbE MAC
 *
 * The implementation is very lightweight. It requires that data in be valid
 * for a packet, once started, until the end of the packet.
 *
 */
/*a To do
 *  Optionally pad short packets
 *  Optionally (configurable) insert timestamp in to packet
 *  Capture timestamp on end of preamble (more predictable than SOP)
 *  Timer to count continuously
 *  Module to retard / accelerate nanosecond timestamp using divide-by-N
 */
/*a Includes */
include "types/timer.h"
include "types/axi.h"
include "types/ethernet.h"

/*a Constants
*/
constant integer preamble_length=8; // 7 of 0x55 one of 0xd5

/*a Types */
/*t t_tx_fsm */
typedef fsm {
    tx_fsm_idle         "Waiting for valid data in";
    tx_fsm_preamble     "Outputting preamble";
    tx_fsm_data         "Outputting data, calculating FCS";
    tx_fsm_fcs          "Outputting FCS";
    tx_fsm_ipg          "Waiting for inter-packet gap";
    tx_fsm_aborting     "Data not valid when required - aborting packet";
    tx_fsm_skipping     "Dropping input data until 'last' asserted";
} t_tx_fsm;

/*t t_tx_action */
typedef enum [5] {
    tx_action_none,
    tx_action_sop                "Packet data valid, send SOP",
    tx_action_preamble           "Send preamble",
    tx_action_preamble_end       "Send last byte of preamble",
    tx_action_data               "Send next byte of packet data and update FCS",
    tx_action_last_data_of_word  "Send last byte of current packet data and update FCS",
    tx_action_data_eop           "Send last byte of packet data and update FCS",
    tx_action_fcs                "Send next byte of FCS",
    tx_action_fcs_end            "Send last byte of FCS",
    tx_action_ipg                "Send idle",
    tx_action_idle               "Start wait for packet data in to be valid",
    tx_action_abort_start        "Send inverted FCS out",
    tx_action_abort              "Send inverted FCS out",
    tx_action_abort_end          "Send inverted FCS out and move to skip",
    tx_action_drop               "Drop any incoming packet data (will not be last)",
    tx_action_drop_idle          "Drop last incoming packet data and move to ipg"
} t_tx_action;

/*t t_fcs_op */
typedef enum [2] {
    fcs_op_none,
    fcs_op_init,
    fcs_op_calc,
    fcs_op_shift
} t_fcs_op;

/*t t_tx_combs */
typedef struct {
    t_tx_action action;
    bit consuming_axi4s;
    bit can_output_symbol;
    bit last_byte_of_packet "Asserted if AXI4S 'last' and last tx strobe";
    bit data_invalid        "Asserted if AXI4S data is not ready for state machine";
    bit[8] axi4s_data_byte;
    bit[8] axi4s_fcs_byte;
    bit[32] next_fcs;
    bit shift_data;
    t_fcs_op fcs_op;
    bit[7] byte_of_packet_plus_one;
} t_tx_combs;

/*t t_tx_state */
typedef struct {
    t_tx_fsm  fsm_state;
    bit[4]    count          "State machine counter";
    t_axi4s32 axi4s          "AXI4S data being consumed";
    t_axi4s32 pending_axi4s  "AXI4S data waiting to be moved to axi4s";
    bit[32]   fcs;
    bit       gmii_tx_valid  "If low, then all GMII TX outputs are low - else to values in gmii_tx";
    t_gmii_tx gmii_tx        "GMII TX data out (if gmii_tx_valid)";
    bit[7]    byte_of_packet "Byte of packet";
    bit[4]    ipg;
} t_tx_state;

/*t t_rx_fsm */
typedef fsm {
    rx_fsm_idle         "Waiting for valid data in";
    rx_fsm_preamble     "Outputting preamble";
    rx_fsm_data         "Outputting data, calculating FCS";
    rx_fsm_wait_for_idle "Waiting for idle from GMII";
} t_rx_fsm;

/*t t_rx_action */
typedef enum [5] {
    rx_action_none,
    rx_action_sop                "Packet data valid, send SOP",
    rx_action_preamble_end       "Send last byte of preamble",
    rx_action_data,
    rx_action_packet_okay,
    rx_action_packet_error,
    rx_action_idle,
    rx_action_overrun,
    rx_action_non_packet_error,
} t_rx_action;

/*t t_rx_combs */
typedef struct {
    t_rx_action action;
    bit[8]  gmii_data;
    bit     gmii_idle;
    bit     gmii_valid_data;
    bit     gmii_valid;
    bit     axi_cannot_take_data;
    bit[32] next_fcs;
    bit fcs_valid;
    bit store_byte;
    bit store_status;
    bit data_ready_for_axi;
    t_fcs_op fcs_op;
    bit[16] byte_of_packet_plus_one;
} t_rx_combs;

/*t t_rx_state */
typedef struct {
    t_axi4s32 axi4s          "AXI4S data being presented";
    t_rx_fsm  fsm_state;
    bit[4] byte_valid;
    bit[32] data_word;
    bit[32]   fcs;
    bit[16]    byte_of_packet "Byte of packet";
    bit[16]    max_mtu        "Largest packet size supported";
} t_rx_state;

/*a Module
*/
/*m gbe_axi4s32 */
module gbe_axi4s32( clock tx_aclk   "Transmit clock domain - AXI-4-S and GMII TX clock",
                    input bit tx_areset_n,
                    input t_axi4s32 tx_axi4s,
                    output bit      tx_axi4s_tready,
                    input   bit gmii_tx_enable "Clock enable for tx_aclk for GMII",
                    output  t_gmii_tx gmii_tx,

                    clock rx_aclk    "Receive clock domain - AXI-4-S and GMII RX clock",
                    input bit rx_areset_n,
                    output t_axi4s32 rx_axi4s,
                    input bit        rx_axi4s_tready,
                    input   bit gmii_rx_enable "Clock enable for rx_aclk for GMII",
                    input   t_gmii_rx gmii_rx,
                    input t_timer_control tx_timer_control "Timer control in TX clock domain"
    )
/*b Documentation */
"""
A light-weight full-duplex Ethernet MAC supporting GMII.

0x04C11DB7  /2= 2608edb /2= 130476d  /2= 9823b6
>>> bits_of_n(32,0x04C11DB7)
[1, 1, 1, 0, 1, 1, 0, 1, 1, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0]
>>> x=bits_of_n(32,0x04C11DB7)
>>> x.reverse()
>>> "%x"%(int_of_bits(x))
0xedb88320 /2= 76dc4190 /2= 3b6e20c8 /2= 1db71064
>>>
                    C704DD7B (bit reverse debb20e3)
7BDD04C7 

"""
/*b Module body */
{
    /*b Tx combs and state */
    comb     t_tx_combs tx_combs;
    clocked clock tx_aclk reset active_low tx_areset_n t_tx_state tx_state = {*=0};

    /*b Tx AXI-4S interface */
    tx_axi4s : {
        tx_axi4s_tready = 1;
        if (tx_combs.shift_data) {
            tx_state.axi4s.t.data[24;0] <= tx_state.axi4s.t.data[24;8];
            tx_state.axi4s.t.strb <= tx_state.axi4s.t.strb>>1;
        }
        if (tx_combs.consuming_axi4s) {
            tx_state.axi4s.valid <= 0;                
        }
        if (tx_state.pending_axi4s.valid) {
            tx_axi4s_tready = 0;
            if (!tx_state.axi4s.valid || tx_combs.consuming_axi4s) {
                tx_state.axi4s               <= tx_state.pending_axi4s;
                tx_state.pending_axi4s.valid <= 0;                
            }
        } elsif (tx_axi4s.valid) {
            tx_state.pending_axi4s <= tx_axi4s;
        }
    }

    /*b Tx state machine */
    tx_fsm : {
        /*b Decode AXI state for FSM */
        tx_combs.data_invalid    = !tx_state.axi4s.valid;
        tx_combs.last_byte_of_packet = (tx_state.axi4s.t.strb<2) && tx_state.axi4s.t.last;
        tx_state.ipg <= 12;
        tx_combs.can_output_symbol = (!tx_state.gmii_tx_valid) || gmii_tx_enable;
        
        /*b TX FSM */
        tx_combs.action = tx_action_none;
        full_switch (tx_state.fsm_state) {
        case tx_fsm_idle: {
            if (tx_state.axi4s.valid && tx_combs.can_output_symbol) {
                tx_combs.action = tx_action_sop;
            }
        }
        case tx_fsm_preamble: {
            if (tx_combs.can_output_symbol) {
                tx_combs.action = tx_action_preamble;
                if (tx_state.count==0) {
                    tx_combs.action = tx_action_preamble_end;
                }
            }
        }
        case tx_fsm_data: {
            if (tx_combs.can_output_symbol) {
                tx_combs.action = tx_action_data;
                if (tx_state.count==0) {
                    tx_combs.action = tx_action_last_data_of_word;
                }
                if (tx_combs.last_byte_of_packet) {
                    tx_combs.action = tx_action_data_eop;
                }
                if (tx_combs.data_invalid) {
                    tx_combs.action = tx_action_abort_start;
                }
            }
        }
        case tx_fsm_fcs: {
            if (tx_combs.can_output_symbol) {
                tx_combs.action = tx_action_fcs;
                if (tx_state.count==0) {
                    tx_combs.action = tx_action_fcs_end;
                }
            }
        }
        case tx_fsm_ipg: {
            if (tx_combs.can_output_symbol) {
                tx_combs.action = tx_action_ipg;
                if (tx_state.count==0) {
                    tx_combs.action = tx_action_idle;
                }
            }
        }
        case tx_fsm_aborting: {
            if (tx_combs.can_output_symbol) {
                tx_combs.action = tx_action_abort;
                if (tx_state.count==0) {
                    tx_combs.action = tx_action_abort_end;
                }
            }
        }
        case tx_fsm_skipping: {
            if (tx_state.axi4s.valid) {
                tx_combs.action = tx_action_drop;
                if (tx_state.axi4s.t.last) {
                    tx_combs.action = tx_action_drop_idle;
                }
            }
        }
        }

        /*b Decode action to state update and other controls
         */
        tx_combs.consuming_axi4s = 0;
        tx_combs.shift_data      = 0;
        tx_combs.fcs_op          = fcs_op_none;
        tx_state.count <= tx_state.count - 1;
        tx_combs.byte_of_packet_plus_one = tx_state.byte_of_packet+1;
        if (tx_state.byte_of_packet==-1) { // Saturate 
            tx_combs.byte_of_packet_plus_one = -1;
        }

        tx_combs.axi4s_data_byte = tx_state.axi4s.t.data[8;0];
        tx_combs.axi4s_data_byte = tx_state.axi4s.t.data[8;0];
        tx_combs.axi4s_fcs_byte  = ~tx_state.fcs[8;0]; 
        if (gmii_tx_enable) {
            tx_state.gmii_tx_valid <= 0;
        }
        
        full_switch (tx_combs.action) {
        case tx_action_none: {
            tx_state.fsm_state <= tx_state.fsm_state;
            tx_state.count     <= tx_state.count;
        }
        case tx_action_sop: {
            tx_state.fsm_state <= tx_fsm_preamble;
            tx_state.gmii_tx_valid <= 1;
            tx_state.gmii_tx.tx_en <= 1;
            tx_state.gmii_tx.tx_er <= 0;
            tx_state.gmii_tx.txd   <= 0x55;
            tx_state.count         <= preamble_length-2; // Since SOP is one, and last preamble byte is different
            tx_state.byte_of_packet <= 0;
            tx_combs.fcs_op         = fcs_op_init;
        }
        case tx_action_preamble: {
            tx_state.gmii_tx_valid <= 1;
        }
        case tx_action_preamble_end: {
            tx_state.fsm_state <= tx_fsm_data;
            tx_state.gmii_tx_valid <= 1;
            tx_state.gmii_tx.txd   <= 0xd5;
            tx_state.count         <= 3;
        }
        case tx_action_data: {
            tx_state.gmii_tx_valid <= 1;
            tx_state.gmii_tx.txd   <= tx_combs.axi4s_data_byte;
            tx_state.byte_of_packet <= tx_combs.byte_of_packet_plus_one;
            tx_combs.shift_data    = 1;
            tx_combs.fcs_op        = fcs_op_calc;
        }
        case tx_action_last_data_of_word: {
            tx_state.gmii_tx_valid <= 1;
            tx_state.gmii_tx.txd   <= tx_combs.axi4s_data_byte;
            tx_state.count         <= 3;
            tx_state.byte_of_packet <= tx_combs.byte_of_packet_plus_one;
            tx_combs.fcs_op        = fcs_op_calc;
            tx_combs.consuming_axi4s = 1;
        }
        case tx_action_data_eop: {
            tx_state.fsm_state <= tx_fsm_fcs;
            tx_state.gmii_tx_valid <= 1;
            tx_state.gmii_tx.txd   <= tx_combs.axi4s_data_byte;
            tx_state.byte_of_packet <= tx_combs.byte_of_packet_plus_one;
            tx_state.count         <= 3;
            tx_combs.fcs_op        = fcs_op_calc;
            tx_combs.consuming_axi4s = 1;
        }
        case tx_action_fcs: {
            tx_state.gmii_tx_valid <= 1;
            tx_state.gmii_tx.txd   <= tx_combs.axi4s_fcs_byte;
            tx_combs.fcs_op        = fcs_op_shift;
        }
        case tx_action_fcs_end: {
            tx_state.fsm_state     <= tx_fsm_ipg;
            tx_state.gmii_tx_valid <= 1;
            tx_state.gmii_tx.txd   <= tx_combs.axi4s_fcs_byte;
            tx_state.count         <= tx_state.ipg;
        }
        case tx_action_ipg: {
            tx_state.fsm_state     <= tx_fsm_ipg;
            tx_state.gmii_tx_valid <= 0;
        }
        case tx_action_idle: {
            tx_state.fsm_state     <= tx_fsm_idle;
            tx_state.gmii_tx_valid <= 0;
        }
        case tx_action_abort_start: {
            tx_state.fsm_state <= tx_fsm_aborting;
            tx_state.count         <= 3;
            tx_state.gmii_tx_valid <= 1;
            tx_state.gmii_tx.txd   <= ~tx_combs.axi4s_fcs_byte;
        }
        case tx_action_abort: {
            tx_state.gmii_tx_valid <= 1;
            tx_state.gmii_tx.txd   <= ~tx_combs.axi4s_fcs_byte;
        }
        case tx_action_abort_end: {
            tx_state.fsm_state <= tx_fsm_skipping;
            tx_state.gmii_tx_valid <= 1;
            tx_state.gmii_tx.txd   <= ~tx_combs.axi4s_fcs_byte;
        }
        case tx_action_drop: {
            tx_state.gmii_tx_valid <= 0;
            tx_combs.consuming_axi4s = 1;
        }
        case tx_action_drop_idle: {
            tx_state.fsm_state <= tx_fsm_ipg;
            tx_state.gmii_tx_valid <= 0;
            tx_combs.consuming_axi4s = 1;
        }
        }

        /*b GMII TX output */
        gmii_tx = {*=0};
        if (tx_state.gmii_tx_valid) {
            gmii_tx = tx_state.gmii_tx;
        }
    }        

    /*b Tx FCS */
    tx_fcs:{
        tx_combs.next_fcs = tx_state.fcs >> 8;
        if (tx_state.fcs[7] ^ tx_combs.axi4s_data_byte[7]) { tx_combs.next_fcs = tx_combs.next_fcs ^ 32hedb88320; }
        if (tx_state.fcs[6] ^ tx_combs.axi4s_data_byte[6]) { tx_combs.next_fcs = tx_combs.next_fcs ^ 32h76dc4190; }
        if (tx_state.fcs[5] ^ tx_combs.axi4s_data_byte[5]) { tx_combs.next_fcs = tx_combs.next_fcs ^ 32h3b6e20c8; }
        if (tx_state.fcs[4] ^ tx_combs.axi4s_data_byte[4]) { tx_combs.next_fcs = tx_combs.next_fcs ^ 32h1db71064; }
        if (tx_state.fcs[3] ^ tx_combs.axi4s_data_byte[3]) { tx_combs.next_fcs = tx_combs.next_fcs ^ 32h0edb8832; }
        if (tx_state.fcs[2] ^ tx_combs.axi4s_data_byte[2]) { tx_combs.next_fcs = tx_combs.next_fcs ^ 32h076dc419; }
        if (tx_state.fcs[1] ^ tx_combs.axi4s_data_byte[1]) { tx_combs.next_fcs = tx_combs.next_fcs ^ 32hee0e612c; }
        if (tx_state.fcs[0] ^ tx_combs.axi4s_data_byte[0]) { tx_combs.next_fcs = tx_combs.next_fcs ^ 32h77073096; }

        full_switch (tx_combs.fcs_op) {
        case fcs_op_init:  { tx_state.fcs <= -1; }
        case fcs_op_calc:  { tx_state.fcs <= tx_combs.next_fcs; }
        case fcs_op_shift: { tx_state.fcs[24;0] <= tx_state.fcs[24;8]; }
        default:           { tx_state.fcs <= tx_state.fcs; }
        }
    }

    /*b Rx combs and state */
    comb     t_rx_combs rx_combs;
    clocked clock rx_aclk reset active_low rx_areset_n t_rx_state rx_state = {*=0};
    /*b Rx state machine */
    rx_fsm : {
        /*b Decode AXI state for FSM */
        rx_combs.gmii_data       = gmii_rx.rxd;
        rx_combs.gmii_idle       = gmii_rx_enable && !gmii_rx.rx_dv && !gmii_rx.rx_er;
        rx_combs.gmii_valid_data = gmii_rx_enable && gmii_rx.rx_dv && !gmii_rx.rx_er;
        rx_combs.gmii_valid      = gmii_rx_enable;

        rx_combs.data_ready_for_axi = 0;
        rx_combs.axi_cannot_take_data = 0;
        if ((rx_state.byte_of_packet[2;0]==0) && rx_state.byte_valid[0]) {
            rx_combs.data_ready_for_axi = 1;
        }
        if (rx_combs.data_ready_for_axi && rx_state.axi4s.valid) {
            rx_combs.axi_cannot_take_data = 1;
        }
        
        /*b RX FSM */
        rx_combs.action = rx_action_none;
        full_switch (rx_state.fsm_state) {
        case rx_fsm_idle: {
            if (rx_combs.gmii_valid_data && (rx_combs.gmii_data==0x55)) {
                rx_combs.action = rx_action_sop;
            } elsif (rx_combs.gmii_valid) {
                rx_combs.action = rx_action_non_packet_error;
            }
        }
        case rx_fsm_preamble: {
            if (rx_combs.gmii_valid_data && (rx_combs.gmii_data==0x55)) {
                rx_combs.action = rx_action_sop;
            } elsif (rx_combs.gmii_valid_data && (rx_combs.gmii_data==0xd5)) {
                rx_combs.action = rx_action_preamble_end;
            } elsif (rx_combs.gmii_valid) {
                rx_combs.action = rx_action_non_packet_error;
            }
        }
        case rx_fsm_data: {
            if (rx_combs.gmii_valid_data) { // rv_dv and not rv_er
                rx_combs.action = rx_action_data;
                if (rx_combs.axi_cannot_take_data) {
                    rx_combs.action = rx_action_overrun;
                }
                if (rx_state.byte_of_packet > rx_state.max_mtu) {
                    rx_combs.action = rx_action_packet_error;
                }
            } elsif (rx_combs.gmii_idle) { // not rx_dv and not rx_er
                rx_combs.action = rx_action_packet_okay; // done without needing more data
                if (rx_combs.fcs_valid) {
                    rx_combs.action = rx_action_packet_error;
                }
            } elsif (rx_combs.gmii_valid) { // rx_er
                rx_combs.action = rx_action_packet_error;
            }
        }
        case rx_fsm_wait_for_idle: {
            if (rx_combs.gmii_idle) {
                rx_combs.action = rx_action_idle;
            }
        }
        }

        /*b Decode action to state update and other controls
         */
        rx_combs.fcs_op          = fcs_op_none;
        rx_combs.byte_of_packet_plus_one = rx_state.byte_of_packet+1;
        rx_combs.store_byte    = 0;
        rx_combs.store_status  = 0;

        full_switch (rx_combs.action) {
        case rx_action_none: {
            rx_state.fsm_state <= rx_state.fsm_state;
        }
        case rx_action_sop: {
            rx_state.fsm_state <= rx_fsm_preamble;
            rx_state.byte_of_packet <= 0;
        }
        case rx_action_preamble_end: {
            rx_state.fsm_state      <= rx_fsm_data;
            rx_state.byte_of_packet <= 0;
            rx_combs.fcs_op          = fcs_op_init;
        }
        case rx_action_data: {
            rx_state.byte_of_packet <= rx_combs.byte_of_packet_plus_one;
            rx_combs.store_byte    = 1;
            rx_combs.fcs_op        = fcs_op_calc;
        }
        case rx_action_packet_okay: { // Packet completed
            rx_state.fsm_state   <= rx_fsm_idle;
            rx_combs.store_status  = 1;
        }
        case rx_action_packet_error: { // Packet completed
            rx_state.fsm_state   <= rx_fsm_wait_for_idle;
            rx_combs.store_status  = 1;
        }
        case rx_action_non_packet_error: { // Packet completed
            rx_state.fsm_state   <= rx_fsm_wait_for_idle;
        }
        case rx_action_idle: { // Packet completed
            rx_state.fsm_state   <= rx_fsm_idle;
        }
        }

        /*b Store data */
        if (rx_state.axi4s.valid && rx_axi4s_tready) {
            rx_state.axi4s.valid <= 0;            
        }
        if (rx_combs.store_byte && rx_combs.data_ready_for_axi) {
            rx_state.axi4s.valid  <= 1;
            rx_state.axi4s.t <= {*=0};
            rx_state.axi4s.t.data <= rx_state.data_word;
            rx_state.axi4s.t.strb <= rx_state.byte_valid;
            rx_state.byte_valid <= 0;
        }
        if (rx_combs.store_byte) {
            full_switch (rx_state.byte_of_packet[2;0]) {
            case 0: {
                rx_state.data_word[8; 0] <= rx_combs.gmii_data;
                rx_state.byte_valid[0]   <= 1;
            }
            case 1: {
                rx_state.data_word[8; 8] <= rx_combs.gmii_data;
                rx_state.byte_valid[1]   <= 1;
            }
            case 2: {
                rx_state.data_word[8;16] <= rx_combs.gmii_data;
                rx_state.byte_valid[2]   <= 1;
            }
            case 3: {
                rx_state.data_word[8;24] <= rx_combs.gmii_data;
                rx_state.byte_valid[3]   <= 1;
            }
            }
        }
        
        /*b GMII RX output */
        rx_axi4s = rx_state.axi4s;
    }        

    /*b Rx FCS */
    rx_fcs:{
        rx_combs.next_fcs = rx_state.fcs >> 8;
        if (rx_state.fcs[7] ^ rx_combs.gmii_data[7]) { rx_combs.next_fcs = rx_combs.next_fcs ^ 32hedb88320; }
        if (rx_state.fcs[6] ^ rx_combs.gmii_data[6]) { rx_combs.next_fcs = rx_combs.next_fcs ^ 32h76dc4190; }
        if (rx_state.fcs[5] ^ rx_combs.gmii_data[5]) { rx_combs.next_fcs = rx_combs.next_fcs ^ 32h3b6e20c8; }
        if (rx_state.fcs[4] ^ rx_combs.gmii_data[4]) { rx_combs.next_fcs = rx_combs.next_fcs ^ 32h1db71064; }
        if (rx_state.fcs[3] ^ rx_combs.gmii_data[3]) { rx_combs.next_fcs = rx_combs.next_fcs ^ 32h0edb8832; }
        if (rx_state.fcs[2] ^ rx_combs.gmii_data[2]) { rx_combs.next_fcs = rx_combs.next_fcs ^ 32h076dc419; }
        if (rx_state.fcs[1] ^ rx_combs.gmii_data[1]) { rx_combs.next_fcs = rx_combs.next_fcs ^ 32hee0e612c; }
        if (rx_state.fcs[0] ^ rx_combs.gmii_data[0]) { rx_combs.next_fcs = rx_combs.next_fcs ^ 32h77073096; }

        full_switch (rx_combs.fcs_op) {
        case fcs_op_init:  { rx_state.fcs <= -1; }
        case fcs_op_calc:  { rx_state.fcs <= rx_combs.next_fcs; }
        default:           { rx_state.fcs <= rx_state.fcs; }
        }
        rx_combs.fcs_valid = (rx_state.fcs==0xdebb20e3); // reverse of 0xC704DD7B 
        rx_state.max_mtu <= -1;
    }

    /*b All done */
}

