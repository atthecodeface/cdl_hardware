/** @copyright (C) 2018,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   tb_riscv_jtag_debug.cdl
 * @brief  Testbench for RISC-V debug over JTAG
 *
 */

/*a Includes
 */
include "jtag.h"
include "apb.h"
include "riscv.h"

/*a External modules */
extern module se_test_harness( clock clk, output t_jtag jtag, output bit tck_enable, input bit tdo )
{
    timing from rising clock clk jtag, tck_enable;
    timing to rising clock clk tdo;
}

typedef struct {
    bit running;
    bit halting;
    bit resuming;
    bit resumed;
    bit attention;
    bit[8] counter;
} t_test_state;

/*a Module
 */
module tb_riscv_jtag_debug( clock jtag_tck,
                          clock apb_clock,
                          input bit reset_n
)
{

    /*b Nets
     */
    net t_jtag jtag;
    net bit tdo;
    net bit[5]ir;
    net t_jtag_action dr_action;
    net bit[50]dr_in;
    net bit[50]dr_tdi_mask;
    net bit[50]dr_out;
    net bit tck_enable;
    comb bit tck_enable_fix;
    gated_clock clock jtag_tck active_high tck_enable_fix jtag_tck_gated;
    net t_riscv_debug_mst debug_mst "Debug master to PDMs";
    clocked clock apb_clock reset active_low reset_n t_riscv_debug_tgt debug_tgt={*=0} "Debug target from PDMs";
    clocked clock apb_clock reset active_low reset_n t_test_state test_state={*=0};

    net  t_apb_request  apb_request  "APB request";
    net t_apb_response apb_response "APB response";

    /*b Instantiate APB timer
     */
    dut_instance: {
        debug_tgt <= {*=0};
        if (debug_mst.valid && (debug_mst.select==0)) {
            debug_tgt <= {valid=1, selected=0, halted=!test_state.running, resumed=test_state.resumed, op_was_none=1};
            test_state.attention <= 0;
        }
        if (test_state.attention) {
            debug_tgt.attention <= 1;
        }
        if (test_state.counter==0) {
            if (test_state.halting) {
                test_state.running <= 0;
                test_state.halting <= 0;
                test_state.attention <= 1;
            }
            if (test_state.resuming) {
                test_state.running <= 1;
                test_state.resuming <= 0;
                test_state.resumed <= 1;
                test_state.attention <= 1;
            }
        } else {
            test_state.counter <= test_state.counter-1;
        }
        if (debug_mst.valid &&(debug_mst.op==rv_debug_set_requests)) {
            test_state.halting <= debug_mst.arg[0];
            test_state.resuming <= debug_mst.arg[1];
            if (!debug_mst.arg[1]) {
                test_state.resumed <= 0;
                test_state.attention <= 1;
            }
            test_state.counter <= 8;
        }
        tck_enable_fix = tck_enable;
        se_test_harness th(clk <- jtag_tck, jtag=>jtag, tck_enable=>tck_enable, tdo<=tdo);

        jtag_tap tap( jtag_tck <- jtag_tck_gated,
                      reset_n <= reset_n,
                      jtag <= jtag,
                      tdo => tdo,

                      ir => ir,
                      dr_action => dr_action,
                      dr_in => dr_in,
                      dr_tdi_mask <= dr_tdi_mask,
                      dr_out <= dr_out );

        riscv_jtag_apb_dm dm_apb( jtag_tck <- jtag_tck_gated,
                      reset_n <= reset_n,

                      ir <= ir,
                      dr_action <= dr_action,
                      dr_in <= dr_in,
                      dr_tdi_mask => dr_tdi_mask,
                      dr_out => dr_out,

                      apb_clock <- apb_clock,
                      apb_request => apb_request,
                      apb_response <= apb_response );

        riscv_i32_debug dm( clk <- apb_clock,
                            reset_n <= reset_n,

                            apb_request <= apb_request,
                            apb_response => apb_response,

                            debug_mst  => debug_mst,
                            debug_tgt <= debug_tgt 
            );
    }
}
