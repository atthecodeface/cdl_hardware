/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   tb_riscv_minimal.cdl
 * @brief  Testbench for minimal RISC-V
 *
 */

/*a Includes
 */
include "srams.h"
include "cpu/riscv/riscv.h"
include "cpu/riscv/riscv_internal_types.h"
include "cpu/riscv/riscv_submodules.h"

/*a External modules */
extern module se_test_harness( clock clk, output t_riscv_i32_coproc_controls  coproc_controls, input t_riscv_i32_coproc_response coproc_response, output t_riscv_config riscv_config)
{
    timing from rising clock clk coproc_controls, riscv_config;
    timing to   rising clock clk coproc_response;
}

/*a Module
 */
module tb_riscv_i32_muldiv( clock clk,
                         input bit reset_n
)
{

    /*b Nets
     */
    net t_riscv_i32_coproc_controls coproc_controls;
    comb t_riscv_i32_coproc_controls coproc_controls_with_feedback;
    net t_riscv_i32_coproc_response coproc_response;
    net t_riscv_config riscv_config;

    /*b Instantiate RISC-V
     */
    riscv_instance: {
        se_test_harness th( clk <- clk,
                            coproc_controls => coproc_controls,
                            coproc_response <= coproc_response,
                            riscv_config => riscv_config );
        
        coproc_controls_with_feedback = coproc_controls;
        coproc_controls_with_feedback.alu_cannot_start    |= coproc_response.cannot_start;
        coproc_controls_with_feedback.alu_cannot_complete |= coproc_response.cannot_complete;
        coproc_controls_with_feedback.dec_to_alu_blocked  |= coproc_response.cannot_start;
        coproc_controls_with_feedback.dec_to_alu_blocked  |= coproc_response.cannot_complete;
        riscv_i32_muldiv dut(  clk <- clk,
                               reset_n <= reset_n,
                               coproc_controls <= coproc_controls_with_feedback,
                               coproc_response => coproc_response,
                               riscv_config <= riscv_config );
    }
}
