/** @copyright (C) 2019,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   clocking_phase_measure.cdl
 * @brief  A module to control a delay module and synchronizer to determine phase length
 *
 * CDL implementation of a module to control a delay module and synchronizer to determine
 * phase length of a clock signal
 *
 * The clock should have as close to a 50-50 duty cycle as possible
 *
 * The module can be prompted to start a measurement; when it does so it will set the
 * delay module to use a zero delay, and it will run through increasing the delay until
 * it gets a consistent value of a synchronized delayed clock for N cycles.
 *
 * It will record this delay and value, then increase the delay again untilt it gets a consistent
 * inverse value. It will then complete the measurement, and report the difference in cycles
 *
 */
/*a Includes */
include "types/encoding.h"

/*a Constants
*/
constant integer qwidth = 10               "1<<qwidth must be >= 8*eye_data_count_running to stop it overflowing";
constant integer eye_data_count_stabilize = 32 "Number of data_clk ticks to wait for stable data after delay has been updated";
constant integer eye_data_count_running   = ((1<<qwidth)/8)-5;
constant integer delay_width = 9;

/*a Types */
/*t t_disparity - encoded with bit[1] = does not change it
     disparity of 00 illegal if disparity in -ve
     disparity of 01 illegal if disparity in +ve
     disparity out = disparity in ^ !disparity[1]
*/
typedef enum[2] {
    disparity_negative = 2b00,                    
    disparity_positive = 2b01,                    
    disparity_zero     = 2b10
} t_disparity;

/*t t_data_6b
*/
typedef struct {
    bit         can_be_control  "Asserted for encodings of 23, 27, 29, 30 and 28";
    bit         can_be_data     "Asserted if symbol is valid data (but may be control if 23/27/29/30)";
    bit[5]      data            "Decoded data value";
    t_disparity disparity       "Disparity of symbol";
} t_data_6b;

/*t t_data_4b
*/
typedef struct {
    bit         valid     "Asserted if a valid 3B4B symbol";
    bit         is_alt    "Asserted if is alt-7";
    bit invert_if_control_and_disparity_minus;
    bit[3]      data      "Decoded data value";
    t_disparity disparity "Disparity of symbol";
} t_data_4b;

/*a Module
*/
/*m decode_8b10b */
module decode_8b10b( input t_8b10b_symbol symbol,
                     output t_8b10b_dec_data dec_data )
"""
This module decodes an 8B10B symbol, splitting it in to two components, each of
which is separately decoded.
"""
{
    comb bit[9] dec_5b6b;
    comb bit[8] dec_3b4b;
    comb t_data_6b data_6b;
    comb t_data_4b data_4b;

    /*b Decode logic */
    decode : {
        /*b Decode 5B6B symbol */
        // Default is neither data nor control
        dec_5b6b = bundle( 2b00,
                           symbol.symbol[5], symbol.symbol[6], symbol.symbol[7], symbol.symbol[8], symbol.symbol[9],
                           2b00 );
        part_switch (symbol.symbol[6;4]) {
            // Data symbols
        case 6b000101: {dec_5b6b = bundle( 2b11, 5d23 , 2b00 ); }
        case 6b000110: {dec_5b6b = bundle( 2b01, 5d8  , 2b00 ); }
        case 6b000111: {dec_5b6b = bundle( 2b01, 5d7  , 2b00 ); }
        case 6b001001: {dec_5b6b = bundle( 2b11, 5d27 , 2b00 ); }
        case 6b001010: {dec_5b6b = bundle( 2b01, 5d4  , 2b00 ); }
        case 6b001011: {dec_5b6b = bundle( 2b01, 5d20 , 2b10 ); }
        case 6b001100: {dec_5b6b = bundle( 2b01, 5d24 , 2b00 ); }
        case 6b001101: {dec_5b6b = bundle( 2b01, 5d12 , 2b10 ); }
        case 6b001110: {dec_5b6b = bundle( 2b01, 5d28 , 2b10 ); }
        case 6b010001: {dec_5b6b = bundle( 2b11, 5d29 , 2b00 ); }
        case 6b010010: {dec_5b6b = bundle( 2b01, 5d2  , 2b00 ); }
        case 6b010011: {dec_5b6b = bundle( 2b01, 5d18 , 2b10 ); }
        case 6b010100: {dec_5b6b = bundle( 2b01, 5d31 , 2b00 ); }
        case 6b010101: {dec_5b6b = bundle( 2b01, 5d10 , 2b10 ); }
        case 6b010110: {dec_5b6b = bundle( 2b01, 5d26 , 2b10 ); }
        case 6b010111: {dec_5b6b = bundle( 2b01, 5d15 , 2b01 ); }
        case 6b011000: {dec_5b6b = bundle( 2b01, 5d0  , 2b00 ); }
        case 6b011001: {dec_5b6b = bundle( 2b01, 5d6  , 2b10 ); }
        case 6b011010: {dec_5b6b = bundle( 2b01, 5d22 , 2b10 ); }
        case 6b011011: {dec_5b6b = bundle( 2b01, 5d16 , 2b01 ); }
        case 6b011100: {dec_5b6b = bundle( 2b01, 5d14 , 2b10 ); }
        case 6b011101: {dec_5b6b = bundle( 2b01, 5d1  , 2b01 ); }
        case 6b011110: {dec_5b6b = bundle( 2b11, 5d30 , 2b01 ); }
        case 6b100001: {dec_5b6b = bundle( 2b11, 5d30 , 2b00 ); }
        case 6b100010: {dec_5b6b = bundle( 2b01, 5d1  , 2b00 ); }
        case 6b100011: {dec_5b6b = bundle( 2b01, 5d17 , 2b10 ); }
        case 6b100100: {dec_5b6b = bundle( 2b01, 5d16 , 2b00 ); }
        case 6b100101: {dec_5b6b = bundle( 2b01, 5d9  , 2b10 ); }
        case 6b100110: {dec_5b6b = bundle( 2b01, 5d25 , 2b10 ); }
        case 6b100111: {dec_5b6b = bundle( 2b01, 5d0  , 2b01 ); }
        case 6b101000: {dec_5b6b = bundle( 2b01, 5d15 , 2b00 ); }
        case 6b101001: {dec_5b6b = bundle( 2b01, 5d5  , 2b10 ); }
        case 6b101010: {dec_5b6b = bundle( 2b01, 5d21 , 2b10 ); }
        case 6b101011: {dec_5b6b = bundle( 2b01, 5d31 , 2b01 ); }
        case 6b101100: {dec_5b6b = bundle( 2b01, 5d13 , 2b10 ); }
        case 6b101101: {dec_5b6b = bundle( 2b01, 5d2  , 2b01 ); }
        case 6b101110: {dec_5b6b = bundle( 2b11, 5d29 , 2b01 ); }
        case 6b110001: {dec_5b6b = bundle( 2b01, 5d3  , 2b10 ); }
        case 6b110010: {dec_5b6b = bundle( 2b01, 5d19 , 2b10 ); }
        case 6b110011: {dec_5b6b = bundle( 2b01, 5d24 , 2b01 ); }
        case 6b110100: {dec_5b6b = bundle( 2b01, 5d11 , 2b10 ); }
        case 6b110101: {dec_5b6b = bundle( 2b01, 5d4  , 2b01 ); }
        case 6b110110: {dec_5b6b = bundle( 2b11, 5d27 , 2b01 ); }
        case 6b111000: {dec_5b6b = bundle( 2b01, 5d7  , 2b01 ); }
        case 6b111001: {dec_5b6b = bundle( 2b01, 5d8  , 2b01 ); }
        case 6b111010: {dec_5b6b = bundle( 2b11, 5d23 , 2b01 ); }

        case 6b001111 : {dec_5b6b = bundle( 2b10, 5d28, 2b01 ); }
        case 6b110000 : {dec_5b6b = bundle( 2b10, 5d28, 2b00 ); }
        }
        data_6b.can_be_control   = dec_5b6b[8];
        data_6b.can_be_data    = dec_5b6b[7];
        data_6b.data           = dec_5b6b[5;2];
        data_6b.disparity      = dec_5b6b[2;0];
    
        /*b Decode 3B4B symbol */
        // Default is neither data nor control
        dec_3b4b = bundle( 1b0, // invert if control and disparity in -ve
                           1b0, // valid
                           1b0, // is alt
                           symbol.symbol[1], symbol.symbol[2], symbol.symbol[3],
                           2b00 );
        part_switch (symbol.symbol[4;0]) {
            // Data symbols (if not a control)
        case 4b0001: {dec_3b4b = bundle( 3b010, 3d7, 2b00);}
        case 4b0010: {dec_3b4b = bundle( 3b010, 3d4, 2b00);}
        case 4b0011: {dec_3b4b = bundle( 3b010, 3d3, 2b10);}
        case 4b0100: {dec_3b4b = bundle( 3b010, 3d0, 2b00);}
        case 4b0101: {dec_3b4b = bundle( 3b110, 3d2, 2b10);} // invert data if control and disparity in -ve
        case 4b0110: {dec_3b4b = bundle( 3b110, 3d6, 2b10);} // invert data if control and disparity in -ve
        case 4b0111: {dec_3b4b = bundle( 3b011, 3d7, 2b01);}
        case 4b1000: {dec_3b4b = bundle( 3b011, 3d7, 2b00);}
        case 4b1001: {dec_3b4b = bundle( 3b110, 3d1, 2b10);} // invert data if control and disparity in -ve
        case 4b1010: {dec_3b4b = bundle( 3b110, 3d5, 2b10);} // invert data if control and disparity in -ve
        case 4b1011: {dec_3b4b = bundle( 3b010, 3d0, 2b01);}
        case 4b1100: {dec_3b4b = bundle( 3b010, 3d3, 2b10);}
        case 4b1101: {dec_3b4b = bundle( 3b010, 3d4, 2b01);}
        case 4b1110: {dec_3b4b = bundle( 3b010, 3d7, 2b01);}
        }
        data_4b.invert_if_control_and_disparity_minus = dec_3b4b[7];
        data_4b.valid          = dec_3b4b[6];
        data_4b.is_alt         = dec_3b4b[5];
        data_4b.data           = dec_3b4b[3;2];
        data_4b.disparity      = dec_3b4b[2;0];

        /*b Decode 8B10B */
        dec_data.valid = (data_6b.can_be_data || data_6b.can_be_control) | data_4b.valid;
        dec_data.data  = bundle(data_4b.data, data_6b.data);
        // note that data of 1,2,5,6 should be ^7 if control AND disparity in is negative
        if ((data_6b.can_be_control && !data_6b.can_be_data) &&
            (symbol.disparity_positive ^ data_6b.disparity[1]) &&
            (data_4b.invert_if_control_and_disparity_minus)
            ) { // only for K.28 really
            dec_data.data  = bundle(~data_4b.data, data_6b.data);
        }

        // control of 28 is allowed with any 3B4B data - and it is marked as can_be_control only
        // control of 23,27,29,30 are allowed only with 3B4B data of alt 7 - these are marked as can_be_control/data
        dec_data.is_control = 0;
        dec_data.is_data  = data_6b.can_be_data;
        if (data_6b.can_be_control) {
            if (!data_6b.can_be_data || data_4b.is_alt) {
                dec_data.is_control = 1;
                dec_data.is_data    = 0;
            }
        }
    
        dec_data.toggles_disparity = (data_4b.disparity[1] != data_6b.disparity[1]);
        dec_data.illegal_if_disparity_negative = 0;
        dec_data.illegal_if_disparity_positive = 0;
        if (data_6b.disparity == disparity_negative) {
            dec_data.illegal_if_disparity_negative = 1;
        } elsif (data_6b.disparity == disparity_positive) {
            dec_data.illegal_if_disparity_positive = 1;
        } else {
            if (data_4b.disparity == disparity_negative) {
                dec_data.illegal_if_disparity_negative = 1;
            } elsif (data_4b.disparity == disparity_positive) {
                dec_data.illegal_if_disparity_positive = 1;
            }
        }

        /*b All done */
        
    }
    /*b All done */
}
