/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   async_reduce_4_60_r
 * @brief  A valid data shift register crossing clock domains
 *
 * Use of the generic_async_reduce module
 *
 * Needs to be built in CDL with the options:
 *
 *  dc:input_width=4
 *
 *  dc:output_width=60
 *
 *  dc:shift_right=1
 *
 *  rmn:generic_async_reduce=async_reduce_4_60_r
 *
 */
/*a Module */
include "generic_async_reduce.cdl"
