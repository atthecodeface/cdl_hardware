/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   riscv_csrs_minimal.cdl
 * @brief  Control/status registers for a minimal RISC-V implementation
 *
 * This file contains a module that implements the in-CPU CSRs
 * required by a RISC-V implementation.
 */

/*a Includes */
include "cpu/riscv/riscv_internal_types.h"

/*a Constants that can be overridden */
constant integer mimpid = 0;
constant integer misa = 0;
constant integer mvendorid = 0;
constant integer mhartid = 0;
constant integer debug_force_disable=0;

/*a Types */
/*t t_csr_write */
typedef struct {
    bit     enable     "Asserted if a CSR write is in progress";
    bit[32] data       "Write data, dependent on current CSR data potentially";
} t_csr_write;

/*t t_mode_combs */
typedef struct {
    bit d;
    bit m;
    bit s;
    bit u;
} t_mode_combs;

/*a Module */
module riscv_csrs_minimal( clock clk                                   "Free-running clock",
                           input bit reset_n                           "Active low reset",
                           input bit riscv_clk_enable                  "RISC-V clock enable",
                           input t_riscv_irqs          irqs            "Interrupts in to the CPU",
                           input t_riscv_csr_access    csr_access      "RISC-V CSR access, combinatorially decoded",
                           output t_riscv_csr_data     csr_data        "CSR respone (including read data), from the current @a csr_access",
                           input t_riscv_csr_controls  csr_controls    "Control signals to update the CSRs",
                           output t_riscv_csrs_minimal csrs            "CSR values"
    )
"""
This module implements a minimal set of RISC-V CSRs, as per v2.1 (May
2016) of the RISC-V instruction set manual user level ISA and v1.9.1
of the privilege architecture (Nov 2016), with the exception that
MTIME has been removed (as this seems to be the correct thing to do).

The privilege specifcation (v1.10) indicates:

* meip is read-only and is derived from the external irq in to this module

* mtip is read-only, cleared by writing to the memory-mapped timer comparator

* msip is read-write in a memory-mapped register somewhere

Hence the irqs structure must provide these three signals


Minimal CSRs as only machine mode and debug mode are supported.
In debug mode every register access is supported.
In machine mode then every register EXCEPT access to ??? is supported.

Given machine mode is the only mode supported:

* there are no SEI and UEI interrupt pins in to this module

* SEIP and UEIP are not supported

* STIP and UTIP are not supported

* SSIP and USIP are not supported

* mstatus.SIE and mstatus.UIE (and previous versions) are hardwired to 0

* mstatus.SPP and mstatus.UPP are hardwired to 0

The mip (machine interrupt pending register) therefore is:

{20b0, MEIP, 3b0, MTIP, 3b0, MSIP, 3b0}

The mie (machine interrupt enable register) is:

{20b0, MEIE, 3b0, MTIE, 3b0, MSIE, 3b0}


The instruction to the pipeline to request an interrupt (which is only
taken if an instruction is in uncommitted in the execution stage) must be generated using the
execution mode and the interrupt enable bits and the interrupt pending
bits.

Hence the 'take interrupt' is (mip & mie) != 0 && mstatus.MIE && (current mode >= machine mode) && (current mode != debug mode).

The required priority order is:

external interrupts, software interrupts, timer interrupts

If an instruction has been committed then it may trap, and the trap
will occur prior to an interrupt which happens after the commit
point. In this case there will be a trap, and the trapped instruction
will be fetched, and then an interrupt can be taken.

When an interrupt is taken the following occurs:

* MPP <= current execution mode (must be machine mode, as debug mode is not interruptible)

* mstatus.MPIE <= mstatus.MIE

Note that WFI should wait independent of mstatus.MIE for (mip & mie) != 0 (given machine mode only)
In debug mode WFI should be a NOP.

WFI may always be a NOP.


User mode interrupts
--------------------

For user mode interrupts there has to be support for delegating an interrupt to user mode - hence the medeleg and mideleg need support (read/write)

User mode interrupts are disabled if mstatus.uie is clear

When an interrupt/exception is delegated to user mode uepc/ucause/utval/mstatus.upie are set to the address, cause etc and mstatus.uie at the interrupt/exception
mstatus.uie is a bit of mstatus that is CLEARED on a user interrupt/exception, and which is set to mstatus.upie on uret; mstatus.upie is then set

uscratch is a 32-bit register for use in the trap handler (and outside it too, if necessary)

utvec is a user vector base for vectored user interrupts

mstatus.uie and mstatus.upie are visible (and only these 2 bits) in 'ustatus'

On uret, uepc/ucause/utval can be cleared (i.e. they are guaranteed to be invalid outside of a user trap handler). mstatus.uie become mstatus.upie; mstatus.upie is set; pc becomes mstatus.uepc

The following CSRs should therefore be supplied for user mode interrupts: ustatus, uie, utvec, uscratch, uepc, ucause, utval, uip.
"""
{

    /*b State
     */
    default clock clk;
    default reset active_low reset_n;
    gated_clock clock clk active_high riscv_clk_enable riscv_clk;
    default clock riscv_clk;
    clocked t_riscv_csrs_minimal csrs={*=0};
    comb t_csr_write  csr_write;
    comb t_mode_combs ret_combs  "Breakout for xRET";
    comb t_mode_combs trap_combs "Breakout for valid trap to mode";

    /*b CSR read/write
     */
    comb bit[32] mstatus;
    comb bit[32] mtvec;
    comb bit[32] mip;
    comb bit[32] mie;
    comb bit[32] dcsr;
    csr_read_write """
    CSR_ADDR_MSTATUS
    CSR_ADDR_MISA
    CSR_ADDR_MVENDORID
    CSR_ADDR_MARCHID
    CSR_ADDR_MIMPID
    CSR_ADDR_MHARTID
    """: {

        /*b Decode read data and 'illegal_access' for the CSR access */
        csr_data = {*=0};
        csr_data.illegal_access = 1;
        mstatus = bundle(csrs.mstatus.sd,
                         8b0,
                         csrs.mstatus.tsr,
                         csrs.mstatus.tw,
                         csrs.mstatus.tvm,
                         csrs.mstatus.mxr,
                         csrs.mstatus.sum,
                         csrs.mstatus.mprv,
                         csrs.mstatus.xs,
                         csrs.mstatus.fs,
                         csrs.mstatus.mpp,
                         2b0,
                         csrs.mstatus.spp,
                         csrs.mstatus.mpie,
                         1b0,
                         csrs.mstatus.spie,
                         csrs.mstatus.upie,
                         csrs.mstatus.mie,
                         1b0,
                         csrs.mstatus.sie,
                         csrs.mstatus.uie
            );
        mie = bundle(20b0,
                     csrs.mie.meip,
                     1b0,
                     csrs.mie.seip,
                     csrs.mie.ueip,
                     csrs.mie.mtip,
                     1b0,
                     csrs.mie.stip,
                     csrs.mie.utip,
                     csrs.mie.msip,
                     1b0,
                     csrs.mie.ssip,
                     csrs.mie.usip );
        mip = bundle(20b0,
                     csrs.mip.meip,
                     1b0,
                     csrs.mip.seip,
                     csrs.mip.ueip,
                     csrs.mip.mtip,
                     1b0,
                     csrs.mip.stip,
                     csrs.mip.utip,
                     csrs.mip.msip,
                     1b0,
                     csrs.mip.ssip,
                     csrs.mip.usip );
        dcsr = bundle(csrs.dcsr.xdebug_ver,
                      12b0,
                      csrs.dcsr.ebreakm,
                      1b0,
                      csrs.dcsr.ebreaks,
                      csrs.dcsr.ebreaku,
                      csrs.dcsr.stepie,
                      csrs.dcsr.stopcount,
                      csrs.dcsr.stoptime,
                      csrs.dcsr.cause,
                      1b0,
                      csrs.dcsr.mprven,
                      csrs.dcsr.nmip,
                      csrs.dcsr.step,
                      csrs.dcsr.prv );
                     
        mtvec = bundle(csrs.mtvec.base, 1b0, csrs.mtvec.vectored);
        part_switch (csr_access.address) {
        case CSR_ADDR_CYCLE     : { csr_data.illegal_access=0; csr_data.read_data = csrs.cycles[32;0]; }
        case CSR_ADDR_CYCLEH    : { csr_data.illegal_access=0; csr_data.read_data = csrs.cycles[32;32]; }
        case CSR_ADDR_MCYCLE    : { csr_data.illegal_access=0; csr_data.read_data = csrs.cycles[32;0]; }
        case CSR_ADDR_MCYCLEH   : { csr_data.illegal_access=0; csr_data.read_data = csrs.cycles[32;32]; }
        case CSR_ADDR_INSTRET   : { csr_data.illegal_access=0; csr_data.read_data = csrs.instret[32;0]; }
        case CSR_ADDR_INSTRETH  : { csr_data.illegal_access=0; csr_data.read_data = csrs.instret[32;32]; }
        case CSR_ADDR_MINSTRET  : { csr_data.illegal_access=0; csr_data.read_data = csrs.instret[32;0]; }
        case CSR_ADDR_MINSTRETH : { csr_data.illegal_access=0; csr_data.read_data = csrs.instret[32;32]; }
        case CSR_ADDR_TIME      : { csr_data.illegal_access=0; csr_data.read_data = csrs.time[32;0]; }
        case CSR_ADDR_TIMEH     : { csr_data.illegal_access=0; csr_data.read_data = csrs.time[32;32]; }
        case CSR_ADDR_MIMPID    : { csr_data.illegal_access=0; csr_data.read_data = mimpid; }
        case CSR_ADDR_MHARTID   : { csr_data.illegal_access=0; csr_data.read_data = mhartid; }
        case CSR_ADDR_MISA      : { csr_data.illegal_access=0; csr_data.read_data = misa; }
        case CSR_ADDR_MVENDORID : { csr_data.illegal_access=0; csr_data.read_data = mvendorid; }
        case CSR_ADDR_MSTATUS   : { csr_data.illegal_access=0; csr_data.read_data = mstatus; }
        case CSR_ADDR_MSCRATCH  : { csr_data.illegal_access=0; csr_data.read_data = csrs.mscratch; }
        case CSR_ADDR_MEPC      : { csr_data.illegal_access=0; csr_data.read_data = csrs.mepc; }
        case CSR_ADDR_MCAUSE    : { csr_data.illegal_access=0; csr_data.read_data = csrs.mcause; }
        case CSR_ADDR_MTVAL     : { csr_data.illegal_access=0; csr_data.read_data = csrs.mtval; }
        case CSR_ADDR_MTVEC     : { csr_data.illegal_access=0; csr_data.read_data = mtvec; } // can be hardwired to any value, or read/write; tests require read-write
            // basic RISC-V tests require the following to not be illegal to write to
        case CSR_ADDR_MEDELEG   : { csr_data.illegal_access=0; csr_data.read_data = 0; } // must be 0 as only machine mode is supported
        case CSR_ADDR_MIDELEG   : { csr_data.illegal_access=0; csr_data.read_data = 0; } // must be 0 as only machine mode is supported
        case CSR_ADDR_MIE       : { csr_data.illegal_access=0; csr_data.read_data = mie; }
        case CSR_ADDR_MIP       : { csr_data.illegal_access=0; csr_data.read_data = mip; }
        case CSR_ADDR_DEPC      : { csr_data.illegal_access=0; csr_data.read_data = csrs.depc; }
        case CSR_ADDR_DCSR      : { csr_data.illegal_access=0; csr_data.read_data = dcsr; }
        }

        /*b Decode CSR writes */
        csr_write.enable = 0;
        csr_write.data = csr_access.write_data;
        if (!csr_access.access_cancelled) {
            part_switch (csr_access.access) {
                case riscv_csr_access_write: { csr_write.enable=1; }
                case riscv_csr_access_rw:    { csr_write.enable=1; }
                case riscv_csr_access_rs:    { csr_write.enable=1; csr_write.data |= csr_data.read_data; }
                case riscv_csr_access_rc:    { csr_write.enable=1; csr_write.data  = csr_data.read_data &~ csr_access.write_data; }
            }
        }

        /*b All done */
    }

    /*b Break out ret and trap */
    ret_trap_breakout: {
        trap_combs = {*=0};
        if (csr_controls.trap.valid) {
            full_switch (csr_controls.trap.to_mode) {
            case rv_mode_debug:      { trap_combs.d = 1; }
            case rv_mode_machine:    { trap_combs.m = 1; }
            case rv_mode_supervisor: { trap_combs.s = 1; }
            case rv_mode_user:       { trap_combs.u = 1; }
            }
            if (debug_force_disable) { trap_combs.m=1; }
        }
        ret_combs = {*=0};
        if (csr_controls.trap.ret) {
            full_switch (csr_controls.trap.cause) {
            case riscv_trap_cause_ret_dret: { ret_combs.d = 1; }
            case riscv_trap_cause_ret_mret: { ret_combs.m = 1; }
            case riscv_trap_cause_ret_sret: { ret_combs.s = 1; }
            case riscv_trap_cause_ret_uret: { ret_combs.u = 1; }
            }
        }
    }
    
    /*b CSR state update */
    csr_state_update """
    """: {
        /*b Mirror time */
        csrs.time <= irqs.time;
            
        /*b Handle CSR cycle state */
        csrs.cycles[32;0] <= csrs.cycles[32;0] + 1;
        if (csrs.cycles[32;0]==-1) {csrs.cycles[32;32] <= csrs.cycles[32;32]+1;}

        if (csr_write.enable && (csr_access.address==CSR_ADDR_MCYCLE)) {
            csrs.cycles[32;0]    <= csr_write.data;
        }
        if (csr_write.enable && (csr_access.address==CSR_ADDR_MCYCLEH)) {
            csrs.cycles[32;32]    <= csr_write.data;
        }

        /*b Handle instruction retire counter state */
        if (csr_controls.retire) {
            csrs.instret[32;0] <= csrs.instret[32;0] + 1;
            if (csrs.instret[32;0]==-1) {csrs.instret[32;32] <= csrs.instret[32;32]+1;}
        }
        if (csr_write.enable && (csr_access.address==CSR_ADDR_MINSTRET)) {
            csrs.instret[32;0] <= csr_write.data;
        }
        if (csr_write.enable && (csr_access.address==CSR_ADDR_MINSTRETH)) {
            csrs.instret[32;32] <= csr_write.data;
        }

        /*b Handle interrupt pending/enable state */
        csrs.mip.meip <= irqs.meip;
        csrs.mip.mtip <= irqs.mtip;
        csrs.mip.msip <= irqs.msip;
        if (csr_write.enable && (csr_access.address==CSR_ADDR_MIE)) {
            csrs.mie.meip <= csr_write.data[11];
            csrs.mie.mtip <= csr_write.data[7];
            csrs.mie.msip <= csr_write.data[3];
        }

        /*b Handle MSTATUS */
        if (trap_combs.m) {
            csrs.mstatus.mpp  <= 2b11; //rv_mode_machine; // Since this is all that is supported; actually 'current mode'
            csrs.mstatus.mpie <= csrs.mstatus.mie;
            csrs.mstatus.mie  <= 0;
        } else {
            if (ret_combs.m) { // note, should enter mode 'csrs.mstatus.mpp'
                csrs.mstatus.mpp  <= 2b11; //rv_mode_machine;
                csrs.mstatus.mpie <= 1;
                csrs.mstatus.mie  <= csrs.mstatus.mpie;
            }
            if (csr_write.enable && (csr_access.address==CSR_ADDR_MSTATUS)) {
                csrs.mstatus.mpp  <= csr_write.data[2;11];
                csrs.mstatus.mpie <= csr_write.data[7];
                csrs.mstatus.mie  <= csr_write.data[3];
            }
        }

        /*b Handle MEPC state */
        if (csr_write.enable && (csr_access.address==CSR_ADDR_MEPC)) {
            csrs.mepc <= csr_write.data;
        }
        if (trap_combs.m) {
            csrs.mepc <= csr_controls.trap.pc;
        }

        /*b Handle MTVEC state */
        if (csr_write.enable && (csr_access.address==CSR_ADDR_MTVEC)) {
            csrs.mtvec.base     <= csr_write.data[30;2];
            csrs.mtvec.vectored <= csr_write.data[0];
        }

        /*b Handle MTVAL state */
        if (trap_combs.m) {
            csrs.mtval <= csr_controls.trap.value;
        }

        /*b Handle MCAUSE state */
        if (csr_write.enable && (csr_access.address==CSR_ADDR_MCAUSE)) {
            csrs.mcause <= csr_write.data;
        }
        if (trap_combs.m) {
            full_switch (csr_controls.trap.cause) {
            case riscv_trap_cause_instruction_misaligned: { csrs.mcause <= bundle(24b0, riscv_mcause_instruction_misaligned); }
            case riscv_trap_cause_instruction_fault:      { csrs.mcause <= bundle(24b0, riscv_mcause_instruction_fault); }
            case riscv_trap_cause_illegal_instruction:    { csrs.mcause <= bundle(24b0, riscv_mcause_illegal_instruction); }
            case riscv_trap_cause_breakpoint:             { csrs.mcause <= bundle(24b0, riscv_mcause_breakpoint); }
            case riscv_trap_cause_load_misaligned:        { csrs.mcause <= bundle(24b0, riscv_mcause_load_misaligned); }
            case riscv_trap_cause_load_fault:             { csrs.mcause <= bundle(24b0, riscv_mcause_load_fault); }
            case riscv_trap_cause_store_misaligned:       { csrs.mcause <= bundle(24b0, riscv_mcause_store_misaligned); }
            case riscv_trap_cause_store_fault:            { csrs.mcause <= bundle(24b0, riscv_mcause_store_fault); }
            case riscv_trap_cause_uecall:                 { csrs.mcause <= bundle(24b0, riscv_mcause_uecall); }
            case riscv_trap_cause_secall:                 { csrs.mcause <= bundle(24b0, riscv_mcause_secall); }
            case riscv_trap_cause_mecall:                 { csrs.mcause <= bundle(24b0, riscv_mcause_mecall); }
            default:                                      { csrs.mcause <= bundle(1b1, 23b0, 4b0, csr_controls.trap.cause[4;0]); } // interrupts
            }
        }

        /*b Handle MSCRATCH state */
        if (csr_write.enable && (csr_access.address==CSR_ADDR_MSCRATCH)) {
            csrs.mscratch <= csr_write.data;
        }

        /*b Handle DSCRATCH state */
        if (csr_write.enable && (csr_access.address==CSR_ADDR_DSCRATCH0)) {
            csrs.dscratch0 <= csr_write.data;
        }
        if (csr_write.enable && (csr_access.address==CSR_ADDR_DSCRATCH1)) {
            csrs.dscratch1 <= csr_write.data;
        }

        /*b Handle DEPC state */
        if (csr_write.enable && (csr_access.address==CSR_ADDR_DEPC)) {
            csrs.depc <= csr_write.data;
        }
        if (trap_combs.d) {
            csrs.depc <= csr_controls.trap.pc;
        }

        /*b Handle DCSR state */
        if (csr_write.enable && (csr_access.address==CSR_ADDR_DCSR)) {
            csrs.dcsr.ebreakm   <= csr_write.data[15];
            csrs.dcsr.ebreaks   <= csr_write.data[13];
            csrs.dcsr.ebreaku   <= csr_write.data[12];
            csrs.dcsr.stepie    <= csr_write.data[11];
            csrs.dcsr.stopcount <= csr_write.data[10];
            csrs.dcsr.stoptime  <= csr_write.data[9];
            csrs.dcsr.mprven    <= csr_write.data[4];
            csrs.dcsr.step      <= csr_write.data[2];
            csrs.dcsr.prv       <= csr_write.data[2;0];
        }
        if (trap_combs.d) {
            csrs.dcsr.cause <= 0;
            csrs.dcsr.prv   <= csr_controls.exec_mode[2;0];
        }
        csrs.dcsr.xdebug_ver <= 4;

        /*b Kill registers if debug not enabled */
        if (debug_force_disable) {
            csrs.depc <= 0;
            csrs.dscratch0 <= 0;
            csrs.dscratch1 <= 0;
            csrs.dcsr <= {*=0};
        }

        /*b Tie-offs for machine mode only */
        //csrs.mtvec.base[;]  <= 0;
        //csrs.mtvec.vectored <= 0;
        csrs.mstatus.mpp    <= 2b11; // only machine mode supported
        csrs.mstatus.sd     <= 0;
        csrs.mstatus.tsr     <= 0;
        csrs.mstatus.tw     <= 0;
        csrs.mstatus.tvm     <= 0;
        csrs.mstatus.mxr     <= 0;
        csrs.mstatus.sum     <= 0;
        csrs.mstatus.mprv     <= 0;
        csrs.mstatus.xs     <= 0;
        csrs.mstatus.fs     <= 0;
        csrs.mstatus.spp     <= 0;
        csrs.mstatus.spie     <= 0;
        csrs.mstatus.upie     <= 0;
        csrs.mstatus.sie     <= 0;
        csrs.mstatus.uie     <= 0;

        csrs.mip.seip     <= 0; // supervisor external interrupt pending from input pin
        csrs.mip.seip_sw  <= 0; // supervisor external interrupt pending from machine mode write
        csrs.mip.ueip     <= 0; // user external interrupt pending from input pin
        csrs.mip.ueip_sw  <= 0; // user external interrupt pending from machine mode write
        csrs.mip.stip     <= 0; // supervisor timer interrupt pending from machine mode write
        csrs.mip.utip     <= 0; // user timer interrupt pending from machine/supervisor mode write
        csrs.mip.ssip     <= 0; // supervisor software interrupt pending from machine/supervisor mode write
        csrs.mip.usip     <= 0; // user software interrupt pending from machine/supervisor mode write

        csrs.mie.seip     <= 0;
        csrs.mie.ueip     <= 0;
        csrs.mie.stip     <= 0;
        csrs.mie.utip     <= 0;
        csrs.mie.ssip     <= 0;
        csrs.mie.usip     <= 0;

        /*b All done */
    }

    /*b Logging */
    logging """
    """: {
        if (csr_write.enable) {
            if (csr_access.address == CSR_ADDR_DSCRATCH0) {
                log("Scratch debug 0 write",
                    "write_data", csr_access.write_data );
            }
        }
    }
}


