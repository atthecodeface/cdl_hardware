/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   riscv_i32_alu.cdl
 * @brief  ALU for i32 RISC-V implementation
 *
 * CDL implementation of RISC-V i32 ALU based on the RISC-V
 * specification v2.1.
 *
 */

/*a Includes
 */
include "cpu/riscv/riscv_pipeline_types.h"
include "cpu/riscv/riscv_internal_types.h"
include "cpu/riscv/riscv.h"

/*a Constants
 */
constant integer coproc_force_disable=0;
constant integer debug_force_disable=0;

/*a Module
 */
module riscv_i32_pipeline_control_flow( input  t_riscv_pipeline_state        pipeline_state,
                                        input  t_riscv_pipeline_response     pipeline_response,
                                        output t_riscv_pipeline_control      pipeline_control,
                                        input t_riscv_i32_coproc_response    coproc_response,
                                        output  t_riscv_mem_access_req       dmem_access_req,
                                        output  t_riscv_csr_access           csr_access,
                                        output t_riscv_i32_coproc_response   pipeline_coproc_response,
                                        input  t_riscv_config                riscv_config
    )
"""

"""
{
    code : {
        pipeline_control.valid = pipeline_state.valid;
        pipeline_control.fetch_action = pipeline_state.fetch_action;
        pipeline_control.fetch_pc = pipeline_state.fetch_pc;
        pipeline_control.mode = pipeline_state.mode;
        pipeline_control.error = pipeline_state.error;
        pipeline_control.tag = pipeline_state.tag;
        pipeline_control.halt = pipeline_state.halt;
        pipeline_control.interrupt_req = pipeline_state.interrupt_req;
        pipeline_control.interrupt_number = pipeline_state.interrupt_number;
        pipeline_control.ebreak_to_dbg = pipeline_state.ebreak_to_dbg;
        pipeline_control.interrupt_to_mode = pipeline_state.interrupt_to_mode;
        pipeline_control.instruction_data = pipeline_state.instruction_data;
        pipeline_control.instruction_debug = pipeline_state.instruction_debug;
        pipeline_control.async_cancel    = pipeline_response.exec.async_cancel;//cannot_complete;

        pipeline_coproc_response = coproc_response;
        if (coproc_force_disable || riscv_config.coproc_disable) {
            pipeline_coproc_response = {*=0};
        }

        pipeline_control.exec_cannot_start    = pipeline_response.exec.cannot_start || pipeline_coproc_response.cannot_start;
        pipeline_control.exec_cannot_complete = pipeline_control.exec_cannot_start  || pipeline_coproc_response.cannot_complete;
        pipeline_control.exec_committed  = pipeline_response.exec.valid && !pipeline_control.exec_cannot_complete;
        pipeline_control.decode_cannot_complete = pipeline_response.decode.valid && pipeline_response.exec.valid && pipeline_control.exec_cannot_complete;

        dmem_access_req = pipeline_response.exec.dmem_access_req;
        // if (!dmem_exec.exec_committed) { dmem_request.access.valid     = 0; }
        if (!pipeline_control.exec_committed) { dmem_access_req.valid = 0; }

        csr_access = pipeline_response.exec.csr_access;
        if (!pipeline_response.exec.valid || pipeline_response.exec.is_illegal) {
            csr_access.access = riscv_csr_access_none;
        }
        csr_access.access_cancelled =  pipeline_response.exec.async_cancel;

    }
}
