/** @copyright (C) 2016-2019,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   timer.cdl
 * @brief  Standardized 64-bit timer with synchronous control
 *
 * CDL implementation of a standard 64-bit timer using synchronous control.
 *
 */
/*a Includes
 */
include "types/apb.h"
include "types/timer.h"

/*a Types */
/*t t_timer_combs
 *
 */
typedef struct {
    bit[5] fractional_sum    "Result of fractional addition, including fractional_bonus";
    bit[33] lower_sum        "Result of integer part of timer, lower bits, summing with timer integer add and fractional overflow";
    bit[32] upper_sum        "Result of upper timer addition - actually an increment based on result of lower_sum carry";
    bit[4]  fractional_half_adder       "Fractional part of half value of interger/fractional adder";
    bit[8]  integer_half_adder          "Integer part of half value of interger/fractional adder";
    bit[5]  fractional_one_and_half_adder       "1-bit int plus fractional part of 3/2 value of interger/fractional adder";
    bit[8]  integer_one_and_half_adder          "Integer part of 3/2 value of interger/fractional adder";
} t_timer_combs;

/*t t_timer_state
 *
 */
typedef struct {
    bit[8]  bonus_subfraction_step "Counter in range 0..denom-1; compared with numer to determine fractional_bonus";
    bit fractional_bonus           "Carry in to timer fractional bonus adder, depending on numer/denom";
    bit[4]  fraction               "Fraction of timer value, accumulating on each enabled cycle";
    bit[32] timer_lower            "Lower 32-bits of integer timer value";
    bit[32] timer_upper            "Upper 32-bits of integer timer value";
    bit     advance                "Last value of timer_control.advance - used in posedge detection";
    bit     retard                 "Last value of timer_control.retard - used in posedge detection";
    bit     hold_adder             "If asserted, hold current adder value";
    bit[4]  fractional_adder       "Fractional adder to use";
    bit[8]  integer_adder          "Integer adder to use";
} t_timer_state;

/*a Module */
module clock_timer( clock clk             "Timer clock",
              input bit reset_n     "Active low reset",
              input t_timer_control timer_control "Control of the timer", 
              output t_timer_value  timer_value
    )
"""
This is a monotonically increasing 64-bit timer with a standard control interface.

The purpose of the timer is to support a 64-bit global nanosecond
clock that can be used as a 'nanoseconds since' an epoch - for PTP
this would be 1 January 1970 00:00:00 TAI, which is 31 December 1969
23:59:51.999918 UTC. A 64-bit nanosecond timestamp with this epoch
wraps roughly in the year 2106.

The timer has a fractional component to permit, for example, a
'nanosecond' timer that is clocked at, say, 600MHz; in this case the
timer is ticked every 1.666ns, and so an addition in each cycle of
0xa to a 4-bit fractional component and a 1 integer component. The
timer_control has, therfore, a fixed-point adder value with a 4-digit
fractional component.

However, this would actually lead to a timer that would be only 99.61% accurate.

Hence a further subfraction capability is supported; this permits a
further 1/16th of a nanosecond (or whatever the timer unit is) to be
added for M out of every N cycles.

In the case of 600MHz a bonus 1/16th should be added for 2 out of
every 3 cycles. This is set using a bonus_subfraction_numer of 0 and a
bonus_subfraction_denom of 2 (meaning for 2 out of every 3 cycles add
a further 1/16th).

Hence every three cycles the timer will have 0x1.b, 0x1.b, 0x1.a
added to it - hence the timer will have gone up by an integer value of
5ns, which is correct for 3 600MHz clock cycles.

If the control values are tied off to zero then the extra fractional
logic will be optimized out.

Some example values for 1ns timer values:

Clock  | Period    | Adder (Int/fraction) | Subfraction Numer/Denom
-------|-----------|----------------------|------------------------
1GHz   |    1ns    |      1 / 0x0         |    0 / 0
800MHz |  1.25ns   |      1 / 0x4         |    0 / 0
600MHz |  1.66ns   |      1 / 0xa         |    0 / 2

The period should be:

  * subfraction numer/denum=0/x: (Int + fraction/16)

  * subfraction numer/denum=M/N: (Int + (fraction+(N-M)/(N+1))/16) 

In addition a synchronous advance/retard option is provided for.
Each time advance is seen going high (i.e. positive edge of advance)
then on an addition the timer will increment by ?.
Each time retard is seen going high the timer will reduces its increment by ?.

Furthermore, there is a synchronize control. When this is asserted, on the next
clock edge where the clock is loaded with the 64-bit synchronization value.

"""
{
    /*b Clock and reset */
    default clock clk;
    default reset active_low reset_n;

    /*b Timer state */
    clocked t_timer_state timer_state= {*=0} "State of the timer and comparator";
    comb    t_timer_combs timer_combs        "Combinatorial decode of timer state and controls";

    /*b Handle the timer and comparator */
    timer_logic """
    The @a timer value can be reset or it may count on a tick, or it
    may just hold its value.

    The timer update logic adds the integer and fractional increments
    to the timer value, with an optional carry (@a fractional_bonus)
    in that is generated and registered on the previous cycle. This
    bonus is one for @a bonus_subfraction_numer out of @a
    bonus_subfraction_denom.

    """: {
        /*b Support advance and retard */
        timer_combs.fractional_half_adder = timer_control.fractional_adder >> 1;
        timer_combs.fractional_half_adder[3] = timer_control.integer_adder[0];
        timer_combs.fractional_one_and_half_adder = bundle(1b0, timer_combs.fractional_half_adder) + bundle(1b0, timer_control.fractional_adder);
        timer_combs.integer_half_adder          = timer_control.integer_adder >> 1;
        timer_combs.integer_one_and_half_adder  = timer_combs.integer_half_adder + timer_control.integer_adder;
        if (timer_combs.fractional_one_and_half_adder[4]) {
            timer_combs.integer_one_and_half_adder  = timer_combs.integer_half_adder + timer_control.integer_adder + 1;
        }
        
        if (!timer_state.hold_adder || timer_control.reset_counter) {
            timer_state.fractional_adder <= timer_control.fractional_adder;
            timer_state.integer_adder    <= timer_control.integer_adder;
            timer_state.hold_adder <= 1;
        }
        if (timer_control.advance && !timer_state.advance) {
            timer_state.fractional_adder <= timer_combs.fractional_one_and_half_adder[4;0];
            timer_state.integer_adder    <= timer_combs.integer_one_and_half_adder;
            timer_state.hold_adder       <= 0;
        } elsif (timer_control.retard && !timer_state.retard) {
            timer_state.fractional_adder <= timer_combs.fractional_half_adder;
            timer_state.integer_adder    <= timer_combs.integer_half_adder;
            timer_state.hold_adder       <= 0;
        }
        if (timer_control.advance || timer_state.advance) {
            timer_state.advance <= timer_control.advance;
        }
        if (timer_control.retard || timer_state.retard) {
            timer_state.retard <= timer_control.retard;
        }
        
        /*b Tick / reset timer */
        timer_combs.fractional_sum = ( bundle(1b0, timer_state.fraction)    +
                                       bundle(1b0, timer_state.fractional_adder) +
                                       (timer_state.fractional_bonus ? 1: 0)
            );
        timer_combs.lower_sum      = ( bundle(1b0, timer_state.timer_lower) +
                                       bundle(25b0, timer_state.integer_adder) +
                                       (timer_combs.fractional_sum[4]?1:0)
            );
        timer_combs.upper_sum      = timer_state.timer_upper;
        if (timer_combs.lower_sum[32]) {
            timer_combs.upper_sum      = timer_state.timer_upper + 1;
        }
        
        if (timer_control.enable_counter) {
            if (timer_control.bonus_subfraction_denom==0) {
                timer_state.bonus_subfraction_step <= 0;
                timer_state.fractional_bonus       <= 0;
            } else {
                timer_state.bonus_subfraction_step <= timer_state.bonus_subfraction_step + 1;
                if (timer_state.bonus_subfraction_step>=timer_control.bonus_subfraction_denom) {
                    timer_state.bonus_subfraction_step <= 0;
                }
                timer_state.fractional_bonus <= 0;
                if (timer_state.bonus_subfraction_step > timer_control.bonus_subfraction_numer) {
                    timer_state.fractional_bonus <= 1;
                }
            }
            timer_state.fraction    <= timer_combs.fractional_sum[4;0];
            timer_state.timer_lower <= timer_combs.lower_sum[32;0];
            timer_state.timer_upper <= timer_combs.upper_sum;
        }
        if (timer_control.reset_counter) {
            timer_state.bonus_subfraction_step <= 0;
            timer_state.fractional_bonus <= 0;
            timer_state.fraction <= 0;
            timer_state.timer_lower <= 0;
            timer_state.timer_upper <= 0;
        }

        /*b Allow synchronization */
        if (timer_control.synchronize[0]) {
            timer_state.timer_lower  <= timer_control.synchronize_value[32; 0];
            timer_state.fraction     <= 0;
        }
        if (timer_control.synchronize[1]) {
            timer_state.timer_upper  <= timer_control.synchronize_value[32;32];
            timer_state.fraction     <= 0;
        }

        /*b Drive outputs */
        timer_value.value = bundle(timer_state.timer_upper, timer_state.timer_lower);
        timer_value.irq = 0;
        timer_value.locked = 0;
    }

    /*b Done
     */
}

/*a Editor preferences and notes
mode: c ***
c-basic-offset: 4 ***
c-default-style: (quote ((c-mode . "k&r") (c++-mode . "k&r"))) ***
outline-regexp: "/\\\*a\\\|[\t ]*\/\\\*[b-z][\t ]" ***
*/
