/** @copyright (C) 2019,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   tb_8b10b.cdl
 * @brief  Testbench for 8b10b encoder and decoder
 *
 */
/*a Includes */
include "types/encoding.h"
include "networking/encoders.h"

/*a External modules */
extern module se_test_harness( clock clk,
                               output t_8b10b_symbol    dec_symbol,
                               output t_8b10b_enc_data  enc_data,
                               input t_8b10b_dec_data  dec_data,
                               input t_8b10b_symbol    enc_symbol
    )
{
    timing to   rising clock clk dec_data, enc_symbol;
    timing from rising clock clk dec_symbol, enc_data;
}

/*a Module */
module tb_8b10b( clock clk,
                 input bit reset_n
)
{
    /*b Nets */
    default clock clk;
    default reset active_low reset_n;
    net t_8b10b_symbol    dec_symbol;
    net t_8b10b_enc_data  enc_data ;
    net t_8b10b_dec_data  dec_data ;
    net t_8b10b_symbol    enc_symbol;
    clocked t_8b10b_dec_data  dec_data_r   = {*=0} ;
    clocked t_8b10b_symbol    enc_symbol_r = {*=0} ;

    /*b Instantiations */
    instantiations: {
        encode_8b10b enc( enc_data <= enc_data,
                          symbol => enc_symbol );
        decode_8b10b dec( symbol <= dec_symbol,
                          dec_data => dec_data);
        se_test_harness th( clk <- clk,
                            enc_data   => enc_data,
                            dec_symbol => dec_symbol,
                            enc_symbol <= enc_symbol_r,
                            dec_data   <= dec_data_r
            );
        enc_symbol_r <= enc_symbol;
        dec_data_r <= dec_data;
        /*b All done */
    }

    /*b All done */
}

