/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   riscv_minimal.cdl
 * @brief  Minimal RISC-V implementation ported to CDL
 *
 * CDL implementation of minimal RISC-V teaching implementation
 *
 * This is a two-stage pipeline implementation, with instruction fetch
 * of the next PC occuring simultaneously with the decode, register
 * read, ALU, data read/write request, data read memory access, and
 * register update.
 *
 * The instruction memory request, then, becomes valid dependent on
 * the decode of the registered instruction last fetched. For most
 * branches this requires only a small amount of logic, but for
 * jump-and-link-register instructions (which uses the full ALU
 * result) this may take a considerable amount of gates to determine
 * the correct branch target and hence next instruction fetch.  Hence
 * the instruction memory request is valid after a considerable delay
 * from the start of the cycle.
 *
 * The return value from the instruction memory request must be valid
 * before the end of the cycle.
 *
 * Any instruction memory implementation must start its access well
 * after the CPU clock edge, , as the request is valid after the CPU
 * clock edge; the resultant read data delay (from the clock edge)
 * then has to be factored in to determine when the next CPU clock
 * edge can occur. Hence it may be sensible to use a double speed
 * clock (e.g. 'fast_clk') to generate CPU clock edges (every other
 * fast_clk edge) and SRAM access clock edges (for a synchronous
 * memory) on the intervening fast_clk edges.
 *
 * The data memory request becomes valid, again, a fair time after the
 * CPU clock edge, as it requires instruction decode, register fetch,
 * and ALU operation to occur prior to the memory address being valid.
 *
 * The data memory response must be valid (for read data!) in the same
 * CPU cycle, as the returning data has to be rotated to the correct
 * byte lanes and prepared for the register file write.
 *
 * Hence a data memory implementation can be similar to that proposed
 * for the instruction memory - that is, accesses start on a memory
 * clock edge that is in the middle of a CPU clock edge, by using a
 * fast_clk.
 *
 */

/*a Includes
 */
include "cpu/riscv/riscv_internal_types.h"
include "cpu/riscv/riscv.h"
include "cpu/riscv/riscv_submodules.h"

/*a Constants
 */
constant integer INITIAL_PC=0x0;

/*a Types
 */
/*t t_ifetch_combs
 *
 * Combinatorials for the instruction fetch
 */
typedef struct {
    t_riscv_pipeline_control_fetch_action fetch_action;
    bit interrupt_req;
    bit[4] interrupt_number;
} t_ifetch_combs;

/*t t_ifetch_state
 *
 * Combinatorials for the instruction fetch
 */
typedef fsm {
    ifetch_fsm_idle;
    ifetch_fsm_restarting;
    ifetch_fsm_fetching;
} t_ifetch_fsm;
typedef struct {
    t_ifetch_fsm state;
    bit running;
    bit[32]      pc    "PC to start fetching from";
} t_ifetch_state;

/*a Module
 */
module riscv_i32_pipeline_control( clock clk,
                                    input bit reset_n,
                                    input t_riscv_csrs_minimal          csrs,
                                    output t_riscv_pipeline_control     pipeline_control,
                                    input t_riscv_pipeline_response   pipeline_response,
                                    input  t_riscv_fetch_resp          ifetch_resp,
                                    input  t_riscv_config              riscv_config,
                                    input t_riscv_i32_trace           trace
)
{
    default clock clk;
    default reset active_low reset_n;
    comb    t_ifetch_combs         ifetch_combs;
    clocked t_ifetch_state         ifetch_state = {*=0, state=ifetch_fsm_idle};
    /*b Pipeline control
     */
    pipeline_control_logic
    """
    The instruction fetch request derives from the
    decode/execute stage (the instruction address that is required
    next) and presents that to the outside world.

    This request may be for any 16-bit aligned address, and two
    successive 16-bit words from that request must be presented,
    aligned to bit 0.

    If the decode/execute stage is invalid (i.e. it does not have a
    valid instruction to decode) then the current PC is requested.
    """:
    {
        if (!ifetch_state.running) { // AND if run from boot time
            ifetch_state.running <= 1;
            ifetch_state.pc <= INITIAL_PC;
        }

        // handle wfi_mode[] too
        //        machine_mode_int_req = 0;
        ifetch_combs.interrupt_req = 0;
        ifetch_combs.interrupt_number = 0;
        if (csrs.mip.mtip & csrs.mie.mtip) {
           ifetch_combs.interrupt_req    = csrs.mstatus.mie; // and only if not in debug
           ifetch_combs.interrupt_number = 7;
        }
        if (csrs.mip.msip & csrs.mie.msip) {
           ifetch_combs.interrupt_req    = csrs.mstatus.mie; // and only if not in debug
           ifetch_combs.interrupt_number = 3;
        }
        if (csrs.mip.meip & csrs.mie.meip) {
           ifetch_combs.interrupt_req    = csrs.mstatus.mie; // and only if not in debug
           ifetch_combs.interrupt_number = 11;
        }

        ifetch_combs.fetch_action   = rv_pc_fetch_action_continue_fetching;
        full_switch (ifetch_state.state) {
        case ifetch_fsm_idle: {
            if (ifetch_state.running) {
                ifetch_state.state <= ifetch_fsm_restarting;
            }
        }
        case ifetch_fsm_restarting: {
            ifetch_combs.fetch_action   = rv_pc_fetch_action_restart_at_pc;
            if (ifetch_resp.valid) {
                ifetch_state.state <= ifetch_fsm_fetching;
            }
        }
            // on a flush NEXT cycle pipeline_response.exec.pc MUST equal ifetch_req.address
            // it always will with this pipeline
        case ifetch_fsm_fetching: { // present request, decode should be valid, pipeline not empty
            ifetch_combs.fetch_action   = rv_pc_fetch_action_continue_fetching;
        }
        }

        pipeline_control = {*=0};
        pipeline_control.valid        = 1;
        pipeline_control.start_pc     = ifetch_state.pc;
        pipeline_control.fetch_action = ifetch_combs.fetch_action;
        pipeline_control.mode  = rv_mode_machine;
        pipeline_control.interrupt_req     = ifetch_combs.interrupt_req;
        pipeline_control.interrupt_number  = ifetch_combs.interrupt_number;
        pipeline_control.interrupt_to_mode = rv_mode_machine;
    }
}
