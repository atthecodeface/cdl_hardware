/** @copyright (C) 2018,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   apb_master_axi.cdl
 * @brief  AXI target to an APB master interface
 *
 * APB master driven by an AXI target (32-bit address, 64-bit data)
 *
 * Supports aligned 32-bit single length transactions only
 *
 * The AXI target supports 32-bit aligned 32-bit read/writes with full
 * byte enables only.
 * 
 * Other transactions should return a slave error response (but they
 * don't as yet)
 *
 */

/*a Includes
 */
include "types/apb.h"
include "types/axi.h"

/*a Types */
/*t t_axi_wr_fsm */
typedef fsm
{
    axi_wr_idle       {
        axi_wr_get_data
            } "Waiting for an AXI write request";
    axi_wr_get_data   {
        axi_wr_do_apb
            } "Waiting for the write data for the write request";
    axi_wr_do_apb     {
        axi_wr_wait_apb
            } "Presenting APB access (when APB is ready)";
    axi_wr_wait_apb   {
        axi_wr_wait_ack
            } "Waiting for APB access to complete";
    axi_wr_wait_ack   {
        axi_wr_idle
            } "Presenting write response to AXI master";
} t_axi_wr_fsm;

/*t t_axi_wr_state */
typedef struct
{
    t_axi_wr_fsm state "State of the AXI write state machine";
    bit     errored    "Asserted if the AXI request did not match the capabilities of the logic";
    bit[12] id         "@a id field of the AXI write request being handled";
    bit[32] address    "@a address of the AXI write request being handled";
    bit[32] data       "@a data from the AXI write data channel for the AXI write request being handled";
} t_axi_wr_state;

/*t t_axi_rd_fsm */
typedef fsm
{
    axi_rd_idle     {
        axi_rd_do_apb
            } "Waiting for an AXI read requests";
    axi_rd_do_apb{
        axi_rd_wait_apb
            } "Requesting an APB read transaction";
    axi_rd_wait_apb{
        axi_rd_wait_ack
            } "Waiting for APB read transaction to complete";
    axi_rd_wait_ack{
        axi_rd_idle
            } "Presenting AXI read response";
} t_axi_rd_fsm;

/*t t_axi_rd_state */
typedef struct
{
    t_axi_rd_fsm state "State of the AXI read state machine";
    bit     errored    "Asserted if the AXI request did not match the capabilities of the logic";
    bit[12] id         "@a id field of the AXI read request being handled";
    bit[32] address    "@a address of the AXI read request being handled";
} t_axi_rd_state;

/*a Module
 */
/*m apb_master_axi
 *
 */
module apb_master_axi( clock aclk                    "AXI and APB clock",
                       input bit areset_n            "AXI and APB reset",
                       input t_axi_request ar        "AXI read request from master",
                       output bit arready            "Ready signal for AXI read requests",
                       input t_axi_request aw        "AXI write request from master",
                       output bit awready            "Ready signal for AXI write requests",
                       input t_axi_write_data w      "AXI write data from master",
                       output bit wready             "Ready signal for write data",
                       input bit bready              "Ready signal from master for returning write responses",
                       output t_axi_write_response b "Write response back to master",
                       input bit rready              "Ready signal from master for returning read data and response",
                       output t_axi_read_response r  "Read response back to master",

                       output t_apb_request     apb_request    "APB request out",
                       input t_apb_response     apb_response   "APB response back"
    )
"""
AXI target mapping to an APB master

This is a very simple AXI target that handles a single AXI transaction
at any one time; it converts this into an APB read or write
transaction, whose completion allows the completion of the AXI
transaction.

This module is currently very primitive, and does not checking of
transaction input really.
"""
{
    /*b Default clock and reset */
    default clock aclk;
    default reset active_low areset_n;

    /*b Clocked state for the AXI inputs from the master - we can accept input if these are not valid */
    clocked bit awready = 0;
    clocked bit arready = 0;
    clocked bit wready = 0;
    clocked t_axi_write_response b={*=0};
    clocked t_axi_read_response  r={*=0};
    clocked t_apb_request apb_request={*=0};

    /*b Clocked state for the AXI state machines */
    clocked t_axi_wr_state axi_wr_state={*=0} "State of the AXI write side";
    clocked t_axi_rd_state axi_rd_state={*=0} "State of the AXI read side";

    /*b Clocked state and decode for the APB transaction side */
    clocked bit apb_access_in_progress = 0  "Asserted if an APB access is in progress";
    comb bit apb_access_start_read          "Asserted if an APB read access should start";
    comb bit apb_access_start_write         "Asserted if an APB write access should start";
    comb bit apb_access_completing          "Asserted if an APB access is completing (psel & penable & pready)";

    /*b AXI-side logic
     *
     * Does not yet check:
     *
     * size must be 32
     * strobes must be all 1
     * burst length must be 0
     * lock must be 0
     * cache must be ?
     * prot must be ?
     * qos / region / user ?
     *
     */
    axi_logic """
    The AXI-side logic has two state machines: one handles AXI write
    requests, the other AXI read requests.

    A write request must be paired with write data, and this permits
    the state machine to then generate a request to the APB side to
    perform an APB write transaction; when that completes, the AXI
    write response can be returned.

    A read request permits the state machine to generate a request to
    the APB side to perform an APB read transaction; when that
    completes, the AXI read response can be returned.

    A read request is only presented if the write state machine is
    idle. Hence @a apb_access_start_write and @a apb_access_start_read
    can never be asserted simultaneously.

    """: {
        arready <= 0;
        wready <= 0;
        apb_access_start_read = 0;
        apb_access_start_write = 0;

        /*b AXI write state machine - idle, get data, do_apb, wait_apb, wait_ack
         */
        full_switch (axi_wr_state.state) {
        case axi_wr_idle: {
            if (aw.valid) {
                awready <= 1;
                wready <= 1;
                axi_wr_state.state <= axi_wr_get_data;
                axi_wr_state.errored <= 0;
                axi_wr_state.id <= aw.id;
                axi_wr_state.address <= aw.addr[32;0];
            }
        }
        case axi_wr_get_data: {
            awready <= 0;
            wready <= 1;
            if (w.valid) {
                if (!w.last) {
                    axi_wr_state.errored <= 1; // max of 1 data cycle
                }
                if (w.last) {
                    wready <= 0;
                    axi_wr_state.state <= axi_wr_do_apb;
                    axi_wr_state.data <= w.data[32;0];
                }
            }
        }
        case axi_wr_do_apb: {
            if (!apb_access_in_progress) {
                apb_access_start_write = 1;
                axi_wr_state.state <= axi_wr_wait_apb;
            }
        }
        case axi_wr_wait_apb: {
            if (apb_access_completing) {
                axi_wr_state.state <= axi_wr_wait_ack;
                b <= {*=0};
                b.valid <= 1;
                b.id <= axi_wr_state.id;
                b.resp <= axi_resp_okay;
            }
        }
        case axi_wr_wait_ack: {
            b.valid <= 1;
            if (bready) {
                b.valid <= 0;
                axi_wr_state.state <= axi_wr_idle;
            }
        }
        }

        /*b AXI reads - rd_idle, rd_do_apb, rd_wait_apb, rd_wait_ack
         *
         * An APB read is only requested if the AXI write state machine is
         * in idle. The AXI write state machine will not request and @a apb_access_start_write
         * in that state, hence @a apb_access_start_read is exclusive with @a apb_access_start_write
         *
         */
        full_switch (axi_rd_state.state) {
        case axi_rd_idle: {
            if (ar.valid) {
                arready <= 1;
                axi_rd_state.state <= axi_rd_do_apb;
                axi_rd_state.errored <= 0;
                axi_rd_state.id <= ar.id;
                axi_rd_state.address <= ar.addr[32;0];
            }
        }
        case axi_rd_do_apb: {
            arready <= 0;
            if (axi_wr_state.state == axi_wr_idle) {
                apb_access_start_read = 1; // apb_access_start_write will not be asserted
                axi_rd_state.state <= axi_rd_wait_apb;
            }
        }
        case axi_rd_wait_apb: {
            if (apb_access_completing) {
                axi_rd_state.state <= axi_rd_wait_ack;
                r <= {*=0};
                r.valid <= 1;
                r.id <= axi_rd_state.id;
                r.resp <= axi_resp_okay; // use apb_request.perr
                r.data <= apb_response.prdata;
                r.last <= 1;
            }
        }
        case axi_rd_wait_ack: {
            r.valid <= 1;
            if (rready) {
                r.valid <= 0;
                axi_rd_state.state <= axi_rd_idle;
            }
        }
        }

        /*b All done */
    }

    /*b APB access logic */
    apb_access_logic """
    An APB access starts with a valid request detected, which drives
    out the APB controls with @p psel high, @p penable low.

    If @p psel is high and @p penable is low then an access must have
    started, and the next clock tick _must_ have penable high.

    If @p psel is high and @p penable is high then the access will continue
    if @p pready is low, but it will complete (with valid read data, if a
    read) if @p pready is high.
    """: {
        apb_access_completing = 0;
        if (apb_access_start_read || apb_access_start_write) {
            apb_access_in_progress <= 1;
            if (apb_access_start_write) {
                apb_request <= { psel=1,
                        pwrite = 1,
                        paddr  = axi_wr_state.address,
                        pwdata = axi_wr_state.data };
            } else {
                apb_request <= { psel=1,
                        pwrite = 0,
                        paddr  = axi_rd_state.address };
            }
        }
        if (apb_request.psel) {
            if (!apb_request.penable) {
                apb_request.penable <= 1;
            } elsif (apb_response.pready) {
                apb_access_completing = 1;
                apb_request.penable <= 0;
                apb_request.psel <= 0;
                apb_access_in_progress <= 0;
            }
        }
    }

    /*b All done */
}
