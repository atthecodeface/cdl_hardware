/** @copyright (C) 2016-2020,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   tb_riscv_minimal.cdl
 * @brief  Testbench for minimal RISC-V
 *
 */

/*a Includes
 */
include "srams.h"
include "types/apb.h"
include "apb/apb_targets.h"
include "cpu/riscv/riscv.h"
include "cpu/riscv/riscv_modules.h"
include "cpu/riscv/riscv_pipeline.h"
include "cpu/riscv/riscv_submodules.h"
include "cpu/riscv/chk_riscv.h"

/*a Types */
/*t t_drop_data */
typedef enum[2] {
    drop_data_none,
    drop_data_16,
    drop_data_32,
    drop_data_all
} t_drop_data;

/*t t_sram_request */
typedef struct {
    bit     valid;
    bit     read_not_write;
    bit[32] address;
    bit[4]  byte_enable;
    bit[32] write_data;
} t_sram_request;

/*t t_inst_combs */
typedef struct {
    bit[64] data_before_drop;
    bit[64] data_after_drop;
    bit[4] half_words_valid;
    bit[4] half_words_will_be_valid;
    t_sram_request sram_request;
    bit request_initial_half;
    t_drop_data drop_data;
} t_inst_combs;

/*t t_inst_state */
typedef struct {
    bit[4]  half_words_valid_before_reading;
    bit     sram_reading;
    bit     initial_half;
    bit[32] address;
    bit[64] data;
} t_inst_state;

/*t t_data_combs */
typedef struct {
    t_sram_request sram_request;
    bit apb_request_valid;
} t_data_combs;

/*t t_data_state */
typedef struct {
    t_riscv_mem_access_req dmem_access_in_progress;
    t_apb_request apb;
} t_data_state;

/*t t_arbiter_combs */
typedef struct {
    t_sram_request sram_request;
    bit grant_to_inst;
    bit grant_to_data;
} t_arbiter_combs;

/*a Module
 */
module riscv_i32_minimal3( clock clk,
                           input bit reset_n,
                           input bit proc_reset_n,
                           input t_riscv_irqs       irqs               "Interrupts in to the CPU",
                           input  t_sram_access_req       sram_access_req,
                           output t_sram_access_resp      sram_access_resp,
                           output t_apb_request           apb_request,
                           input  t_apb_response          apb_response,
                           input  t_riscv_debug_mst       debug_mst,
                           output t_riscv_debug_tgt       debug_tgt,
                           input  t_riscv_config          riscv_config,
                           output t_riscv_i32_trace       trace
)
"""
An instantiation of Reve-R with multiplier coprocessor and debug, with a single SRAM

Compressed instructions are supported IF i32c_force_disable is 0 and riscv_config.i32c is 1
Multiply/divide coprocesor is supported IF i32c_force_disable is 0 and riscv_config.i32m is 1

A single memory is used for instruction and data, at address 0

Any access outside of the bottom 1MB is passed as a request out of this module.
"""
{
    /*b Default clock and reset
     */
    default clock clk;
    default reset active_low reset_n;

    /*b Nets
     */
    net   t_riscv_debug_tgt debug_tgt;
    net   t_riscv_i32_trace       trace;

    net  t_riscv_mem_access_req  dmem_access_req;
    comb t_riscv_mem_access_resp dmem_access_resp;

    net  t_riscv_fetch_req  rv_imem_access_req;
    comb t_riscv_fetch_resp rv_imem_access_resp;
    net t_riscv_csr_controls      csr_controls;
    net t_riscv_csr_data          csr_data;
    net t_riscv_csr_access        csr_access;
    net t_riscv_csrs              csrs;

    /*b Nets for the pipeline
     */
    net t_riscv_pipeline_state        pipeline_state;
    net t_riscv_pipeline_control      pipeline_control;
    net t_riscv_pipeline_response     pipeline_response;
    net t_riscv_pipeline_fetch_req    pipeline_fetch_req;
    net t_riscv_pipeline_fetch_data   pipeline_fetch_data;
    net t_riscv_pipeline_trap_request pipeline_trap_request;

    /*b State and comb
     */
    comb    t_inst_combs inst_combs;
    clocked t_inst_state inst_state = {*=0};
    comb    t_data_combs data_combs;
    clocked t_data_state data_state = {*=0};
    comb    t_arbiter_combs arbiter_combs;
    net bit[32] sram_read_data;

    net t_riscv_i32_coproc_controls  coproc_controls;
    net t_riscv_i32_coproc_response  coproc_response;
    net t_riscv_i32_coproc_response  pipeline_coproc_response;

    /*b SRAM and arbiter */
    sram_and_arbiter: {
        arbiter_combs.grant_to_inst = 0;
        arbiter_combs.grant_to_data = 0;

        arbiter_combs.sram_request = data_combs.sram_request;
        if (data_combs.sram_request.valid) {
            arbiter_combs.grant_to_data = 1;
            arbiter_combs.sram_request  = data_combs.sram_request;
        } elsif (inst_combs.sram_request.valid) {
            arbiter_combs.grant_to_inst = 1;
            arbiter_combs.sram_request = inst_combs.sram_request;
        } else {
            arbiter_combs.sram_request.valid = 0;
        }
        sram_access_resp = {*=0};

        /*b SRAM instance */
        se_sram_srw_16384x32_we8 mem(sram_clock     <- clk,
                                     select         <= arbiter_combs.sram_request.valid,
                                     read_not_write <= arbiter_combs.sram_request.read_not_write,
                                     write_enable   <= arbiter_combs.sram_request.byte_enable,
                                     address        <= arbiter_combs.sram_request.address[14;2],
                                     write_data     <= arbiter_combs.sram_request.write_data,
                                     data_out       => sram_read_data );
    }

    /*b Instruction memory
     */
    srams: {
        /*b Create data buffer value from SRAM read data and current valid data buffer */
        inst_combs.data_before_drop = inst_state.data;
        inst_combs.half_words_valid = inst_state.half_words_valid_before_reading;
        if (inst_state.sram_reading) {
            inst_combs.half_words_valid = inst_state.half_words_valid_before_reading + 2;
            if    (inst_state.half_words_valid_before_reading==0) { inst_combs.data_before_drop[32;0]  = sram_read_data; }
            elsif (inst_state.half_words_valid_before_reading==1) { inst_combs.data_before_drop[32;16] = sram_read_data; }
            else                                                  { inst_combs.data_before_drop[32;32] = sram_read_data; }
            assert (inst_state.half_words_valid_before_reading<=2, "Incorrect value for half_words_valid_before_reading if we are reading");
            if (inst_state.initial_half) {
                inst_combs.data_before_drop[16;0] = sram_read_data[16;16];
                inst_combs.half_words_valid = 1;
            }
        }

        /*b Decode amount of data to drop given request */
        inst_combs.drop_data = drop_data_none;
        full_switch (rv_imem_access_req.req_type) {
        case rv_fetch_none: {
            inst_combs.drop_data = drop_data_all;
        }
        case rv_fetch_nonsequential: {
            inst_combs.drop_data = drop_data_all;
        }
        case rv_fetch_repeat: {
            inst_combs.drop_data = drop_data_none;
        }
        case rv_fetch_sequential_16: {
            inst_combs.drop_data = drop_data_16;
        }
        case rv_fetch_sequential_32: {
            inst_combs.drop_data = drop_data_32;
        }
        }

        /*b Decode amount of data valid after drop */
        inst_combs.half_words_will_be_valid = inst_combs.half_words_valid;
        inst_combs.data_after_drop          = inst_combs.data_before_drop;
        full_switch (inst_combs.drop_data) {
        case drop_data_none: {
            inst_combs.half_words_will_be_valid = inst_combs.half_words_valid;
        }
        case drop_data_16: {
            inst_combs.data_after_drop[48;0] = inst_combs.data_before_drop[48;16];
            if    (inst_combs.half_words_valid==0) { inst_combs.half_words_will_be_valid = 0; }
            elsif (inst_combs.half_words_valid==1) { inst_combs.half_words_will_be_valid = 0; }
            elsif (inst_combs.half_words_valid==2) { inst_combs.half_words_will_be_valid = 1; }
            elsif (inst_combs.half_words_valid==3) { inst_combs.half_words_will_be_valid = 2; }
            else                                   { inst_combs.half_words_will_be_valid = 3; }
        }
        case drop_data_32: {
            inst_combs.data_after_drop[32;0] = inst_combs.data_before_drop[32;32];
            if    (inst_combs.half_words_valid==0) { inst_combs.half_words_will_be_valid = 0; }
            elsif (inst_combs.half_words_valid==1) { inst_combs.half_words_will_be_valid = 0; }
            elsif (inst_combs.half_words_valid==2) { inst_combs.half_words_will_be_valid = 0; }
            elsif (inst_combs.half_words_valid==3) { inst_combs.half_words_will_be_valid = 1; }
            else                                   { inst_combs.half_words_will_be_valid = 2; }
        }
        case drop_data_all: {
            inst_combs.half_words_will_be_valid = 0;
        }
        }

        /*b Decode address to fetch and whether it is valid */
        inst_combs.sram_request = {*=0};
        inst_combs.request_initial_half = 0;
        inst_combs.sram_request.read_not_write  = 1;
        inst_combs.sram_request.address         = inst_state.address;
        full_switch (rv_imem_access_req.req_type) {
        case rv_fetch_none: {
            inst_combs.sram_request.valid = 0;
            inst_combs.request_initial_half  = 0;
        }
        case rv_fetch_nonsequential: {
            inst_combs.sram_request.valid        = 1;
            inst_combs.request_initial_half      = rv_imem_access_req.address[1];
            inst_combs.sram_request.address      = rv_imem_access_req.address;
        }
        default: {
            inst_combs.request_initial_half   = inst_state.initial_half;
            inst_combs.sram_request.valid     = (inst_combs.half_words_will_be_valid<=2);
            inst_combs.sram_request.address   = inst_state.address;
            if (inst_state.sram_reading) {
                inst_combs.request_initial_half   = 0;
                inst_combs.sram_request.address   = inst_state.address+4;
            }
        }
        }

        /*b Present response */
        rv_imem_access_resp          = {*=0};
        rv_imem_access_resp.data     = inst_combs.data_after_drop[32;0];
        if (rv_imem_access_req.req_type!=rv_fetch_none) {
            if (inst_combs.half_words_will_be_valid>=2) {
                rv_imem_access_resp.valid = 1;
            }
        }

        /*b Update state */
        inst_state.data                            <= inst_combs.data_after_drop;
        inst_state.sram_reading                    <= arbiter_combs.grant_to_inst && inst_combs.sram_request.valid;
        inst_state.initial_half                    <= inst_combs.request_initial_half;
        inst_state.half_words_valid_before_reading <= inst_combs.half_words_will_be_valid;
        inst_state.address                         <= inst_combs.sram_request.address;

    }

    /*b Data memory
     */
    data_memory: {
        /*b Decode data request */
        data_combs.apb_request_valid       = 0;
        data_combs.sram_request.valid      = 0;
        data_combs.sram_request.read_not_write = (dmem_access_req.req_type != rv_mem_access_write);
        data_combs.sram_request.address        = dmem_access_req.address;
        data_combs.sram_request.byte_enable    = dmem_access_req.byte_enable;
        data_combs.sram_request.write_data     = dmem_access_req.write_data;
        if (dmem_access_req.valid) {
            data_combs.sram_request.valid          = 1;
            if (dmem_access_req.address[12;20]!=0) { // 3h0xxxxxxx is SRAM, rest is APB
                data_combs.sram_request.valid      = 0;
                data_combs.apb_request_valid       = 1;
            }
        }

        /*b Generate dmem_access_resp and update APB transaction state */
        dmem_access_resp = {*=0};
        dmem_access_resp.ack             = 1;
        dmem_access_resp.access_complete = 1;
        dmem_access_resp.may_still_abort = 0;
        dmem_access_resp.abort_req       = 0;
        dmem_access_resp.read_data       = sram_read_data;
        if (data_state.apb.penable) {
            dmem_access_resp.read_data   = apb_response.prdata;
        }

        if (data_state.apb.psel) {
            dmem_access_resp.ack             = 0;
            dmem_access_resp.access_complete = 0;
            dmem_access_resp.may_still_abort = 1;
            data_state.apb.penable <= 1;
            if (data_state.apb.penable) {
                dmem_access_resp.abort_req = apb_response.perr;
                if (apb_response.pready || apb_response.perr) {
                    dmem_access_resp.ack             = 1;
                    dmem_access_resp.access_complete = 1;
                }
            }
        }

        /*b Update state */
        data_state.dmem_access_in_progress.valid <= 0;
        if (dmem_access_resp.ack) {
            data_state.apb.psel    <= 0;
            data_state.apb.penable <= 0;
            if (dmem_access_req.valid) {
                data_state.dmem_access_in_progress <= dmem_access_req;
                if (data_combs.apb_request_valid) {
                    data_state.apb.psel    <= 1;
                    data_state.apb.pwrite  <= (dmem_access_req.req_type == rv_mem_access_write);
                    data_state.apb.pwdata  <= dmem_access_req.write_data;
                    data_state.apb.paddr   <= dmem_access_req.address;
                }
            }
        }

        /*b APB request out */
        apb_request = data_state.apb;

        /*b All done */
    }

    /*b Instantiate Reve-R pipeline
     */
    reve_r_pipeline: {
        riscv_i32_pipeline_control pc(clk       <- clk,
                                      riscv_clk <- clk,
                                      reset_n          <= reset_n,
                                      riscv_clk_enable <= 1,
                                      csrs <= csrs,
                                      pipeline_state => pipeline_state,
                                      pipeline_response <= pipeline_response,
                                      pipeline_fetch_data <= pipeline_fetch_data,
                                      pipeline_control <= pipeline_control,
                                      riscv_config     <= riscv_config,
                                      trace            <= trace,
                                      debug_mst        <= debug_mst,
                                      debug_tgt        => debug_tgt,
                                      rv_select <= 0 );

        riscv_i32_pipeline_control_fetch_req pc_fetch_req( pipeline_state <= pipeline_state,
                                                           pipeline_response <= pipeline_response,
                                                           pipeline_fetch_req => pipeline_fetch_req,
                                                           ifetch_req => rv_imem_access_req );

        riscv_i32_pipeline_control_fetch_data pc_fetch_data( pipeline_state <= pipeline_state,
                                                             ifetch_req  <= rv_imem_access_req,
                                                             ifetch_resp <= rv_imem_access_resp,
                                                             pipeline_fetch_req <= pipeline_fetch_req,
                                                             pipeline_fetch_data => pipeline_fetch_data );

        riscv_i32_pipeline_trap_interposer ti( pipeline_state         <= pipeline_state,
                                               pipeline_response      <= pipeline_response,
                                               dmem_access_resp       <= dmem_access_resp,
                                               pipeline_trap_request  => pipeline_trap_request,
                                               riscv_config           <= riscv_config
        );

        riscv_i32_pipeline_control_flow cf( pipeline_state <= pipeline_state,
                                            ifetch_req  <= rv_imem_access_req,
                                            pipeline_response <= pipeline_response,
                                            pipeline_trap_request  <= pipeline_trap_request,
                                            coproc_response <= coproc_response,
                                            pipeline_control => pipeline_control,
                                            dmem_access_resp <= dmem_access_resp,
                                            dmem_access_req => dmem_access_req,
                                            csr_access     => csr_access,
                                            pipeline_coproc_response => pipeline_coproc_response,
                                            coproc_controls  => coproc_controls,
                                            csr_controls     => csr_controls,
                                            trace            => trace,
                                            riscv_config <= riscv_config
        );

        riscv_i32c_pipeline3 pipe( clk <- clk,
                                  reset_n <= reset_n,
                                  pipeline_control <= pipeline_control,
                                  pipeline_response => pipeline_response,
                                  pipeline_fetch_data <= pipeline_fetch_data,
                                  dmem_access_resp <= dmem_access_resp,
                                  coproc_response <= pipeline_coproc_response,
                                  csr_read_data    <= csr_data.read_data,
                                  riscv_config <= riscv_config);

    }

    /*b CSRs
     */
    csr_instance: {
        riscv_csrs_machine_debug_user_irq csrs( clk       <- clk,
                                                riscv_clk <- clk,
                                                reset_n <= reset_n,
                                                riscv_clk_enable <= 1,
                                                irqs <= irqs,
                                                csr_access     <= csr_access,
                                                csr_data       => csr_data,
                                                csr_controls   <= csr_controls,
                                                csrs => csrs
            );
    }

    /*b Coprocessors
     */
    coprocessors: {
        riscv_i32_muldiv m( clk <- clk,
                            reset_n <= reset_n,
                            coproc_controls <= coproc_controls,
                            coproc_response => coproc_response,
                            riscv_config <= riscv_config );

    }

    /*b Checkers - for matching trace etc
     */
    checkers: {
        chk_riscv_ifetch checker_ifetch( clk <- clk,
                                         fetch_req <= rv_imem_access_req,
                                         fetch_resp <= rv_imem_access_resp
                                         //error_detected =>,
                                         //cycle => ,
            );
        chk_riscv_trace checker_trace( clk <- clk,
                                       trace <= trace
                                         //error_detected =>,
                                         //cycle => ,
            );
    }

    /*b All done
     */
}
