/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   riscv_minimal.cdl
 * @brief  Minimal RISC-V implementation ported to CDL
 *
 * CDL implementation of minimal RISC-V teaching implementation
 *
 * This is a two-stage pipeline implementation, with instruction fetch
 * of the next PC occuring simultaneously with the decode, register
 * read, ALU, data read/write request, data read memory access, and
 * register update.
 *
 * The instruction memory request, then, becomes valid dependent on
 * the decode of the registered instruction last fetched. For most
 * branches this requires only a small amount of logic, but for
 * jump-and-link-register instructions (which uses the full ALU
 * result) this may take a considerable amount of gates to determine
 * the correct branch target and hence next instruction fetch.  Hence
 * the instruction memory request is valid after a considerable delay
 * from the start of the cycle.
 *
 * The return value from the instruction memory request must be valid
 * before the end of the cycle.
 *
 * Any instruction memory implementation must start its access well
 * after the CPU clock edge, , as the request is valid after the CPU
 * clock edge; the resultant read data delay (from the clock edge)
 * then has to be factored in to determine when the next CPU clock
 * edge can occur. Hence it may be sensible to use a double speed
 * clock (e.g. 'fast_clk') to generate CPU clock edges (every other
 * fast_clk edge) and SRAM access clock edges (for a synchronous
 * memory) on the intervening fast_clk edges.
 *
 * The data memory request becomes valid, again, a fair time after the
 * CPU clock edge, as it requires instruction decode, register fetch,
 * and ALU operation to occur prior to the memory address being valid.
 *
 * The data memory response must be valid (for read data!) in the same
 * CPU cycle, as the returning data has to be rotated to the correct
 * byte lanes and prepared for the register file write.
 *
 * Hence a data memory implementation can be similar to that proposed
 * for the instruction memory - that is, accesses start on a memory
 * clock edge that is in the middle of a CPU clock edge, by using a
 * fast_clk.
 *
 */

/*a Includes
 */
include "riscv.h"
include "riscv_modules.h"
include "srams.h"

/*a Types
 */
/*t t_riscv_clock_phase
 *
 * Phase of the RISC-V clock, dependent on the imem/dmem requests it performs
 */
typedef fsm {
    rcp_clock_high          "RISC-V clock high; decode of instruction presents correct dmem/imem requests for the whole RISC-V cycle";
    rcp_dread_in_progress   "RISC-V clock low with data memory read in progress; will do instruction fetch next";
    rcp_dwrite_in_progress  "RISC-V clock low with data memory write in progress; will do instruction fetch next or clock will go high";
    rcp_ifetch_in_progress  "RISC-V clock low with fetch of instruction, clock will go high";
    rcp_clock_low           "RISC-V clock low with no requests from RISC-V, will go high";
} t_riscv_clock_phase;

/*t t_ifetch_src */
typedef enum[2] {
    ifetch_src_sram,
    ifetch_src_reg
} t_ifetch_src;

/*t t_data_src */
typedef enum[2] {
    data_src_sram,
    data_src_reg,
    data_src_access
} t_data_src;

/*t t_riscv_clock_action
 */
typedef enum[3] {
    riscv_clock_action_rise,
    riscv_clock_action_fall,
    riscv_clock_action_ifetch,
    riscv_clock_action_dread,
    riscv_clock_action_dwrite,
    riscv_clock_action_wait
} t_riscv_clock_action;

/*a Module
 */
module riscv_i32_minimal( clock clk,
                          input bit reset_n,
                          input t_riscv_irqs       irqs               "Interrupts in to the CPU",
                          output t_riscv_mem_access_req  data_access_req,
                          input  t_riscv_mem_access_resp data_access_resp,
                          input  t_sram_access_req       sram_access_req,
                          output t_sram_access_resp      sram_access_resp,
                          input  t_riscv_config          riscv_config,
                          output t_riscv_i32_trace       trace
)
"""
An instantiation of the single stage pipeline RISC-V with RV32I with a single SRAM

Compressed instructions are not supported

A single memory is used for instruction and data, at address 0

Any access outside of the bottom 1MB is passed as a request out of this module.
"""
{

    /*b State and comb
     */
    default clock clk;
    default reset active_low reset_n;

    net t_riscv_fetch_req       ifetch_req;
    comb  t_riscv_fetch_resp    ifetch_resp;
    net t_riscv_i32_trace       trace_pipe;
    net t_riscv_i32_coproc_controls  coproc_controls;
    comb t_riscv_i32_coproc_response   coproc_response;
    comb  t_riscv_config          riscv_config_pipe;
    net  t_riscv_mem_access_req  dmem_access_req;
    comb t_riscv_mem_access_resp dmem_access_resp;
    clocked bit[32] ifetch_reg = 0;

    comb  t_riscv_mem_access_req  data_sram_access_req;
    clocked t_riscv_mem_access_req  data_access_req = {*=0};

    comb t_riscv_mem_access_req  imem_access_req;
    comb t_riscv_mem_access_resp imem_access_resp;

    /*b State and comb
     */
    net bit[32] mem_read_data;
    comb t_riscv_mem_access_req   mem_access_req;
    comb t_ifetch_src ifetch_src;
    comb t_data_src data_src;
    comb bit sram_access_ack;
    clocked t_sram_access_req  sram_access_req_r = {*=0};
    clocked t_sram_access_resp sram_access_resp = {*=0};

    /*b Clock control
     */
    comb bit riscv_clk_enable;
    clocked t_riscv_clock_phase riscv_clock_phase=rcp_clock_high;
    comb t_riscv_clock_action riscv_clock_action;
    clocked clock clk reset active_low reset_n bit riscv_clk_high = 0;
    gated_clock clock clk active_high riscv_clk_enable riscv_clk;
    clock_control """
    The clock control for a single SRAM implementation could be
    performed with three high speed clocks for each RISC-V
    clock. However, this is a slightly more sophisticated design.

    A minimal RISC-V clock cycle requires at most one instruction fetch and at
    most one of data read or data write.

    With a synchronous memory, a memory read must be presented to the
    SRAM at high speed clock cycle n-1 if the data is to be valid at
    the end of high speed clock cycle n.

    So if just an instruction fetch is required then a first high
    speed cycle is used to present the ifetch, and a second high speed
    cycle is the instruction being read. This is presented directly to
    the RISC-V core.

    If an instruction fetch and data read are required then a first
    high speed cycle is used to present the data read, a second to
    present the ifetch and perform the data read - with the data out
    registered at the start of a third high speed cycle while the
    instruction being read. This is presented directly to the RISC-V
    core; the data read is presented from its stored register

    To ease implementation, and because the minimal RISC-V probably
    always requests an instruction fetch, if a data fetch only is
    requested then the flow follows as if an instruction fetch had
    been requested.

    If an instruction fetch and data write are required then a
    first high speed cycle is used to present the data write, a second
    to present the ifetch and perform the data write, and a third high
    speed cycle while the instruction being read. This is presented
    directly to the RISC-V core.
    """ : {
        data_sram_access_req = dmem_access_req;
        if (dmem_access_req.address[12;20]!=0) {
            data_sram_access_req.read_enable = 0;
            data_sram_access_req.write_enable = 0;
        }
        if (riscv_clk_high) { // first cycle of riscv_clk
            data_access_req.read_enable <= 0;
            data_access_req.write_enable <= 0;
            if (dmem_access_req.read_enable || dmem_access_req.write_enable) {
                data_access_req <= dmem_access_req;
            }
            if (dmem_access_req.address[12;20]==0) {
                data_access_req.read_enable <= 0;
                data_access_req.write_enable <= 0;
            }
        } else {
            if (data_access_req.read_enable || data_access_req.write_enable) {
                if (!data_access_resp.wait) {
                    data_access_req.read_enable <= 0;
                    data_access_req.write_enable <= 0;
                }
            }
        }

        riscv_clock_action = riscv_clock_action_rise;
        ifetch_src = ifetch_src_sram;
        data_src   = data_src_access;
        full_switch (riscv_clock_phase) {
        case rcp_clock_high: { // riscv_clk has just gone high, so core is presenting memory requests
            riscv_clock_action = riscv_clock_action_fall; // might be doing a data access ?
            if (imem_access_req.read_enable) {
                riscv_clock_action = riscv_clock_action_ifetch;
            } else {
                if (data_sram_access_req.read_enable) {
                    riscv_clock_action = riscv_clock_action_dread;
                } elsif (data_sram_access_req.write_enable) {
                    riscv_clock_action = riscv_clock_action_dwrite;
                }
            }
        }
        case rcp_clock_low: {
            ifetch_src = ifetch_src_reg;
            riscv_clock_action = riscv_clock_action_rise; // or wait for data access to complete
            if ((data_access_req.read_enable || data_access_req.write_enable) && data_access_resp.wait) {
                riscv_clock_action = riscv_clock_action_wait;
            }
        }
        case rcp_ifetch_in_progress: {
            riscv_clock_action = riscv_clock_action_rise; // or wait for data access to complete
            if ((data_access_req.read_enable || data_access_req.write_enable) && data_access_resp.wait) {
                riscv_clock_action = riscv_clock_action_wait;
            }
            if (data_sram_access_req.read_enable) {
                riscv_clock_action = riscv_clock_action_dread;
            } elsif (data_sram_access_req.write_enable) {
                riscv_clock_action = riscv_clock_action_dwrite;
            }
        }
        case rcp_dwrite_in_progress: {
            riscv_clock_action = riscv_clock_action_rise;
            ifetch_src = ifetch_src_reg;
        }
        case rcp_dread_in_progress: {
            riscv_clock_action = riscv_clock_action_rise;
            ifetch_src = ifetch_src_reg;
            data_src   = data_src_sram;
        }
        }

        riscv_clk_enable = 0;
        full_switch (riscv_clock_action) {
        case riscv_clock_action_fall: {
            riscv_clock_phase <= rcp_clock_low;
        }
        case riscv_clock_action_rise: { 
            riscv_clock_phase <= rcp_clock_high;
            riscv_clk_enable = 1;
        }
        case riscv_clock_action_wait: { 
            riscv_clock_phase <= rcp_clock_low; // it is possibly already low; make sure it is there
        }
        case riscv_clock_action_ifetch: { 
            riscv_clock_phase <= rcp_ifetch_in_progress;
        }
        case riscv_clock_action_dread: { 
            riscv_clock_phase <= rcp_dread_in_progress;
        }
        case riscv_clock_action_dwrite: { 
            riscv_clock_phase <= rcp_dwrite_in_progress;
        }
        }
        riscv_clk_high <= riscv_clk_enable;
    }

    /*b Instantiate srams
     *
     * SRAM access path can run when no RISC-V access is required.
     *
     * However, RISC-V could run a large number of stores or loads
     * So the SRAM access path can also usurp the dread/dwrite, and potentially hold them off
     *  
     */
    srams: {
        sram_access_ack = 1;
        mem_access_req = {*=0, address=data_sram_access_req.address, byte_enable=data_sram_access_req.byte_enable, write_data=data_sram_access_req.write_data};
        full_switch (riscv_clock_action) {
        case riscv_clock_action_dread: {
            mem_access_req = {read_enable=1, address=data_sram_access_req.address};
        }
        case riscv_clock_action_dwrite: {
            mem_access_req = {write_enable=1, byte_enable=data_sram_access_req.byte_enable, address=data_sram_access_req.address, write_data=data_sram_access_req.write_data};
        }
        case riscv_clock_action_ifetch: {
            mem_access_req = {read_enable=imem_access_req.read_enable, address=imem_access_req.address};
        }
        default: {
            if (sram_access_req_r.valid) {
                mem_access_req = {address=sram_access_req_r.address[32;0], byte_enable=sram_access_req_r.byte_enable[4;0], write_data=sram_access_req_r.write_data[32;0]};
                sram_access_ack = 1;
            }
        }
        }
        se_sram_srw_16384x32_we8 mem(sram_clock <- clk,
                                     select         <= mem_access_req.read_enable || mem_access_req.write_enable,
                                     read_not_write <= mem_access_req.read_enable,
                                     write_enable   <= mem_access_req.write_enable ? mem_access_req.byte_enable:4b0,
                                     address        <= mem_access_req.address[14;2],
                                     write_data     <= mem_access_req.write_data,
                                     data_out       => mem_read_data );
        if (sram_access_resp.ack) {
            sram_access_resp.valid <= 1;
            sram_access_resp.id    <= sram_access_req_r.id;
            sram_access_resp.data[32;0]  <= mem_read_data;
        }
        if (sram_access_req.valid) {
            sram_access_req_r <= sram_access_req;
        }
        if (sram_access_ack) {
            sram_access_req_r.valid <= 0;
        }
        if (sram_access_resp.ack || sram_access_ack) {
            sram_access_resp.ack <= sram_access_ack;
        }
        
        if (riscv_clock_phase==rcp_ifetch_in_progress) {
            ifetch_reg <= mem_read_data;
        }

        imem_access_resp.wait       = 0;
        imem_access_resp.read_data  = mem_read_data;
        if (ifetch_src == ifetch_src_reg) {
            imem_access_resp.read_data  = ifetch_reg;
        }
        dmem_access_resp.wait = 0;
        dmem_access_resp.read_data = data_access_resp.read_data;
        if (data_src == data_src_sram) {
            dmem_access_resp.read_data = mem_read_data;
        }
    }

    /*b Ifetch stage
     */
    instruction_fetch_stage: {
        imem_access_req             = {*=0};
        imem_access_req.read_enable = ifetch_req.valid;
        imem_access_req.address     = bundle(1b0,ifetch_req.address[31;1]);
        imem_access_req.address     = ifetch_req.address;
        ifetch_resp = {*=0};
        ifetch_resp.valid = ifetch_req.valid && !imem_access_resp.wait;
        ifetch_resp.data  = imem_access_resp.read_data;
    }

    /*b Pipeline */
    pipeline: {
        coproc_response = {*=0};
        riscv_config_pipe = riscv_config;
        riscv_config_pipe.i32c = 0;
        riscv_config_pipe.i32m = 0;
        riscv_i32c_pipeline pipeline(clk              <- riscv_clk,
                                     reset_n          <= reset_n,
                                     irqs             <= irqs,
                                     ifetch_req       => ifetch_req,
                                     ifetch_resp      <= ifetch_resp,
                                     dmem_access_req  => dmem_access_req,
                                     dmem_access_resp <= dmem_access_resp,
                                     coproc_controls  => coproc_controls,
                                     coproc_response  <= coproc_response,
                                     riscv_config     <= riscv_config_pipe,
                                     trace            => trace_pipe );
        trace = trace_pipe;
        trace.instr_valid    = trace_pipe.instr_valid    && riscv_clk_enable;
        trace.rfw_data_valid = trace_pipe.rfw_data_valid && riscv_clk_enable;
    }

    /*b All done */
}

