/** @copyright (C) 2019,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   vcu108_riscv.cdl
 * @brief  RISC-V design for the VCU108 board
 *

 */

/*a Includes
 */
include "types/video.h"
include "types/apb.h"
include "types/csr.h"
include "types/dprintf.h"
include "types/sram.h"
include "types/uart.h"
include "types/memories.h"
include "types/subsystem.h"
include "srams.h"
include "apb/apb_targets.h"
include "apb/apb_masters.h"
include "csr/csr_targets.h"
include "csr/csr_masters.h"
include "utils/dprintf_modules.h"
include "utils/async_reduce_modules.h"
include "video/framebuffer_modules.h"

typedef bit[32] t_bit32;
typedef struct {
    bit uart_src_dprintf;
    bit video_src_debug;
} t_debug;

/*a Constants */
constant integer num_dprintf_requesters=8;

/*a Module
 */
/*m subsys_minimal
 *
 * Subsystem with APB modules that can be used as a common block
 *
 */
module subsys_minimal( clock clk,
                       input bit reset_n,

                       input  t_apb_request     master_apb_request "APB request from main system",
                       output t_apb_response    master_apb_response "APB request from main system",
                       input  t_dprintf_req_4   master_dprintf_req "Dprintf request from board (sync to clk)",
                       output bit               master_dprintf_ack "Ack for dprintf request",
                       output t_csr_request     master_csr_request,
                       input  t_csr_response    master_csr_response,

                       input  t_subsys_inputs   subsys_inputs,
                       output t_subsys_outputs  subsys_outputs,

                       clock video_clk,
                       input bit video_reset_n,
                       output t_video_bus video_bus,
                       input bit        tx_axi4s_tready,
                       output t_axi4s32 tx_axi4s,
                       input t_axi4s32  rx_axi4s,
                       output bit       rx_axi4s_tready,
                       output t_timer_control timer_control,
                       input bit[32] analyzer_trace
    )
{
    /*b Clock and reset */
    default clock clk;
    default reset active_low reset_n;

    /*b Nets and combs for APB */
    net t_apb_response master_apb_response;
    net  t_apb_request proc_apb_request;
    net t_apb_response proc_apb_response;
    net  t_apb_request apb_request;

    comb bit[4]        apb_request_sel;
    comb bit           apb_request_apb "Asserted if APB selected and to the local APB";
    comb bit           apb_request_csr "Asserted if APB selected and to the CSR bus";
    comb t_apb_request timer_apb_request;
    comb t_apb_request gpio_apb_request;
    comb t_apb_request i2c_apb_request;
    comb t_apb_request uart_apb_request;
    comb t_apb_request dprintf_apb_request;
    comb t_apb_request csr_apb_request;
    comb t_apb_request fb_sram_apb_request;
    comb t_apb_request dprintf_uart_apb_request;
    comb t_apb_request axi4s_apb_request;
    comb t_apb_request anal_apb_request;

    net t_apb_response  timer_apb_response;
    net t_apb_response  gpio_apb_response;
    net t_apb_response  i2c_apb_response;
    net t_apb_response  uart_apb_response;
    net t_apb_response  dprintf_apb_response;
    net t_apb_response  csr_apb_response;
    net t_apb_response  fb_sram_apb_response;
    net t_apb_response  dprintf_uart_apb_response;
    net t_apb_response  axi4s_apb_response;
    net t_apb_response  anal_apb_response;
    comb t_apb_response apb_response;

    /*b Timer controls etc */
    clocked t_timer_control timer_control={*=0};
    net     t_timer_control rv_timer_control;
    net  t_timer_value timer_value;
    net bit[16] gpio_output;
    net bit[16] gpio_output_enable;
    clocked bit[16]  gpio_input=0;
    net bit     gpio_input_event;
    net bit[32] fb_sram_ctrl;
    clocked t_debug debug={*=0};

    /*b Dprintf requests and muxing */
    net  t_dprintf_req_4 apb_dprintf_req "Dprintf request from APB target";
    comb bit             apb_dprintf_ack "Ack for dprintf request from APB target";

    net bit[num_dprintf_requesters]                 dprintf_ack;
    clocked t_dprintf_req_4[num_dprintf_requesters] dprintf_req={*=0};
    net bit[num_dprintf_requesters-1]               mux_dprintf_ack "Ack for dprintf request after multiplexing";
    net t_dprintf_req_4[num_dprintf_requesters-1]   mux_dprintf_req "Dprintf request after multiplexing";

    net  bit                                        fifo_dprintf_ack_fb   "Ack for dprintf request after multiplexing";
    net  bit                                        fifo_dprintf_ack_uart "Ack for dprintf request after multiplexing";
    comb t_dprintf_req_4                            fifo_dprintf_req_fb   "Dprintf request after multiplexing";
    comb t_dprintf_req_4                            fifo_dprintf_req_uart "Dprintf request after multiplexing";

    comb bit                                        fifo_dprintf_ack "Ack for dprintf request after multiplexing";
    net t_dprintf_req_4                             fifo_dprintf_req "Dprintf request after multiplexing";
    net t_dprintf_byte dprintf_byte;

    net t_csr_request   csr_request;
    comb t_csr_response csr_response;
    clocked t_csr_response csr_response_r = {*=0};
    net t_csr_response tt_debug_framebuffer_csr_response;
    net t_csr_response tt_vga_framebuffer_csr_response;
    net t_csr_response timeout_csr_response;
    comb t_sram_access_req tt_display_sram_access_req;
    net t_video_bus vga_video_bus;
    net t_video_bus debug_video_bus;

    clocked t_apb_processor_request  apb_processor_request={*=0};
    clocked bit                      apb_processor_completed = 0;
    net t_apb_processor_response  apb_processor_response;
    net t_apb_rom_request         apb_rom_request;
    net bit[40]                   apb_rom_data;

    net t_sram_access_req  fb_sram_access_req;
    comb t_sram_access_resp fb_sram_access_resp;

    comb t_uart_rx_data  uart_rx;
    net   t_uart_tx_data uart_tx;
    net   t_uart_status  uart_status;

    net t_i2c i2c_master;

    /*b AXI */
    net bit       rx_axi4s_tready;
    net t_axi4s32 tx_axi4s;

    net  t_sram_access_req  tx_sram_access_req  "SRAM access request";
    net  t_sram_access_req  rx_sram_access_req  "SRAM access request";
    clocked t_sram_access_resp rx_sram_access_resp ={*=0} "SRAM access response";
    net bit[32] rx_sram_read_data;
    clocked t_sram_access_req  rx_current_sram_access={*=0}  "SRAM access request";
    clocked t_sram_access_resp tx_sram_access_resp ={*=0} "SRAM access response";
    net bit[32] tx_sram_read_data;
    clocked t_sram_access_req  tx_current_sram_access={*=0}  "SRAM access request";

    net bit[32] analyzer_mux_control;
    
    /*b APB processor */
    apb_processor_instances: {
        apb_processor_request.address <= 0;
        apb_processor_request.valid   <= !apb_processor_completed;
        if (apb_processor_response.acknowledge) {
            apb_processor_request.valid   <= 0;
            apb_processor_completed <= 1;
        }

        apb_processor apbp( clk <- clk,
                            reset_n <= reset_n,

                            apb_processor_request <= apb_processor_request,
                            apb_processor_response => apb_processor_response,
                            apb_request   => proc_apb_request,
                            apb_response  <= proc_apb_response,
                            rom_request   => apb_rom_request,
                            rom_data      <= apb_rom_data );

        se_sram_srw_256x40 apb_rom(sram_clock <- clk,
                                   select <= apb_rom_request.enable,
                                   address <= apb_rom_request.address[8;0],
                                   read_not_write <= 1,
                                   write_data <= 0,
                                   data_out => apb_rom_data );

    }

    /*b APB master multiplexing and decode */
    apb_multiplexing_decode: {
        apb_master_mux apb_mux_rp( clk <- clk,
                               reset_n <= reset_n,
                               apb_request_0 <= master_apb_request,
                               apb_request_1 <= proc_apb_request,

                               apb_response_0 => master_apb_response,
                               apb_response_1 => proc_apb_response,

                               apb_request =>  apb_request,
                               apb_response <= apb_response );

        apb_request_sel          = apb_request.paddr[4;16]; // 2MB of address space, [4;16] as select
        apb_request_apb          = apb_request.psel && !apb_request.paddr[20];  // 1MB of address space, [20]==0
        apb_request_csr          = apb_request.psel &&  apb_request.paddr[20];   // 1MB of address space, [20]==1
        timer_apb_request        = apb_request;
        gpio_apb_request         = apb_request;
        dprintf_apb_request      = apb_request;
        uart_apb_request         = apb_request;
        fb_sram_apb_request      = apb_request;
        dprintf_uart_apb_request = apb_request;
        i2c_apb_request          = apb_request;
        axi4s_apb_request        = apb_request;
        anal_apb_request         = apb_request;
        csr_apb_request          = apb_request;

        timer_apb_request.paddr        = apb_request.paddr >> 2;
        gpio_apb_request.paddr         = apb_request.paddr >> 2;
        dprintf_apb_request.paddr      = apb_request.paddr >> 2;
        uart_apb_request.paddr         = apb_request.paddr >> 2;
        fb_sram_apb_request.paddr      = apb_request.paddr >> 2;
        dprintf_uart_apb_request.paddr = apb_request.paddr >> 2;
        i2c_apb_request.paddr          = apb_request.paddr >> 2;
        axi4s_apb_request.paddr        = apb_request.paddr >> 2;
        anal_apb_request.paddr         = apb_request.paddr >> 2;

        timer_apb_request.psel        = apb_request_apb && (apb_request_sel==0);
        gpio_apb_request.psel         = apb_request_apb && (apb_request_sel==1);
        dprintf_apb_request.psel      = apb_request_apb && (apb_request_sel==2);
        fb_sram_apb_request.psel      = apb_request_apb && (apb_request_sel==7);
        uart_apb_request.psel         = apb_request_apb && (apb_request_sel==9);
        dprintf_uart_apb_request.psel = apb_request_apb && (apb_request_sel==10);
        i2c_apb_request.psel          = apb_request_apb && (apb_request_sel==12);
        axi4s_apb_request.psel        = apb_request_apb && (apb_request_sel==13);
        anal_apb_request.psel         = apb_request_apb && (apb_request_sel==14);
        
        csr_apb_request.psel          = apb_request_csr;
        csr_apb_request.paddr[16;16]  = bundle(12b0,apb_request.paddr[4;16]);
        csr_apb_request.paddr[16;0]   = bundle( 2b0,apb_request.paddr[14;2]);

        apb_response = {*=0, pready=1};
        apb_response |= timer_apb_response;
        apb_response |= gpio_apb_response;
        apb_response |= uart_apb_response;
        apb_response |= axi4s_apb_response;
        apb_response |= anal_apb_response;
        apb_response |= dprintf_apb_response;
        apb_response |= dprintf_uart_apb_response;
        apb_response |= i2c_apb_response;
        apb_response |= csr_apb_response;
        apb_response.pready = 1;
        apb_response.pready = apb_response.pready & gpio_apb_response.pready;
        apb_response.pready = apb_response.pready & uart_apb_response.pready;
        apb_response.pready = apb_response.pready & axi4s_apb_response.pready;
        apb_response.pready = apb_response.pready & anal_apb_response.pready;
        apb_response.pready = apb_response.pready & dprintf_apb_response.pready;
        apb_response.pready = apb_response.pready & dprintf_uart_apb_response.pready;
        apb_response.pready = apb_response.pready & i2c_apb_response.pready;
        apb_response.pready = apb_response.pready & csr_apb_response.pready;
        if (apb_request_sel==7) { apb_response = fb_sram_apb_response; }
    }

    /*b Dprintf requesting */
    dprintf_requesting : {
        for (i; num_dprintf_requesters) {
            if (dprintf_ack[i]) {
                dprintf_req[i].valid <= 0;
            }
        }

        if (apb_request.psel && apb_request.penable && apb_response.pready) {
            dprintf_req[1] <= {valid=1, address=40,
                    data_0=bundle(40h41_50_42_3a_80, 7b0,apb_request.pwrite, 16h_20_87), // APB:%x %08x %08x %08x (pwrite paddr pwdata prdata)
                    data_1=bundle(apb_request.paddr, 32h20000087),
                    data_2=bundle(apb_request.pwdata, 32h20000087),
                    data_3=bundle(apb_response.prdata,    8hff, 24h0) };
        }
        if (csr_request.valid && csr_response.acknowledge) {
            dprintf_req[2] <= {valid=1, address=80,
                    data_0=bundle(40h43_53_52_3a_80, 7b0,csr_request.read_not_write, 16h_20_83), // CSR:%x %04x %04x %08x (read_not_write select address data)
                    data_1=bundle(csr_request.select,  48h200000000083),
                    data_2=bundle(csr_request.address, 48h200000000087),
                    data_3=bundle(csr_request.data,    8hff, 24h0) };
        }
        if (rx_sram_access_req.valid && rx_sram_access_resp.ack) {
            dprintf_req[3] <= {valid=1, address=120,
                    data_0=bundle(40h52_58_53_3a_81, rx_sram_access_req.id,16h_20_80), // RXS:%x %x %08x %08x %x (id read_not_write address data be)
                    data_1=bundle(7b0,rx_sram_access_req.read_not_write,  56h20000000000087),
                    data_2=bundle(rx_sram_access_req.address,    32h20000087),
                    data_3=bundle(rx_sram_access_req.write_data[32;0], 16h2080, rx_sram_access_req.byte_enable, 8hff) };
        }
        if (rx_sram_access_resp.valid) {
            dprintf_req[4] <= {valid=1, address=160,
                    data_0=bundle(40h52_58_53_3a_81, rx_sram_access_resp.id,16h_20_87), // RXS:%x %x %08x %08x %x (id read_data)
                    data_1=bundle(rx_sram_access_resp.data[32;0], 8hff, 24h0) };
        }

        apb_dprintf_ack = 1;
        if (dprintf_req[0].valid) {
            apb_dprintf_ack = 0;
            if (dprintf_ack[0]) {
                dprintf_req[0].valid <= 0;
            }
        } else {
            if (apb_dprintf_req.valid) {
                dprintf_req[0]  <= apb_dprintf_req;
            }
        }
        
        master_dprintf_ack = 1;
        if (dprintf_req[7].valid) {
            master_dprintf_ack = 0;
            if (dprintf_ack[7]) {
                dprintf_req[7].valid <= 0;
            }
        } else {
            if (master_dprintf_req.valid) {
                dprintf_req[7] <= master_dprintf_req;
            }
        }

        for (i; num_dprintf_requesters) {
            if (fb_sram_ctrl[i] && !subsys_inputs.switches[2]) {
                dprintf_req[i].valid <= 0;
            }
        }

        debug.video_src_debug  <= subsys_inputs.switches[0];
        debug.uart_src_dprintf <= subsys_inputs.switches[1];
        if (fb_sram_ctrl[16]) {
            debug.uart_src_dprintf <= fb_sram_ctrl[17];
        }
        
    }

    /*b Dprintf multiplexing */
    dprintf_multiplexing """
    mux[n-2] = req[n-2] * req[n-1]
    mux[n-3] = req[n-2] * mux[n-2]
    mux[2]   = req[2] * mux[3]
    mux[1]   = req[1] * mux[2]
    mux[0]   = req[0] * mux[1]
    """: {
        dprintf_4_mux tdm_n( clk <- clk,
                             reset_n <= reset_n,
                             req_a <= dprintf_req[num_dprintf_requesters-2],
                             ack_a => dprintf_ack[num_dprintf_requesters-2],
                             req_b <= dprintf_req[num_dprintf_requesters-1],
                             ack_b => dprintf_ack[num_dprintf_requesters-1],
                             req => mux_dprintf_req[num_dprintf_requesters-2],
                             ack <= mux_dprintf_ack[num_dprintf_requesters-2] );

        for (i; num_dprintf_requesters-2) {
            dprintf_4_mux tdm[i]( clk <- clk, reset_n <= reset_n,
                                  req_a <= dprintf_req[i],
                                  ack_a => dprintf_ack[i],
                                  req_b <= mux_dprintf_req[i+1],
                                  ack_b => mux_dprintf_ack[i+1],
                                  req => mux_dprintf_req[i],
                                  ack <= mux_dprintf_ack[i] );
        }
        dprintf_4_fifo_4 dpf( clk <- clk, reset_n <= reset_n,
                            req_in <= mux_dprintf_req[0],
                            ack_in => mux_dprintf_ack[0],
                            req_out => fifo_dprintf_req,
                            ack_out <= fifo_dprintf_ack );

    }

    /*b APB targets */
    apb_target_instances: {
        apb_target_sram_interface fb_sram_if( clk <- clk,
                                           reset_n <= reset_n,
                                           apb_request  <= fb_sram_apb_request,
                                           apb_response => fb_sram_apb_response,
                                           sram_ctrl    => fb_sram_ctrl,
                                           sram_access_req => fb_sram_access_req,
                                           sram_access_resp <= fb_sram_access_resp );

        apb_target_dprintf apb_dprintf( clk <- clk,
                                    reset_n <= reset_n,
                                    apb_request  <= dprintf_apb_request,
                                    apb_response => dprintf_apb_response,
                                    dprintf_req => apb_dprintf_req,
                                    dprintf_ack <= apb_dprintf_ack );

        apb_target_rv_timer timer( clk <- clk,
                                   reset_n <= reset_n,
                                   timer_control <= timer_control,
                                   apb_request  <= timer_apb_request,
                                   apb_response => timer_apb_response,
                                   timer_value => timer_value,
                                    timer_control_out => rv_timer_control );

        apb_target_gpio gpio( clk <- clk,
                              reset_n <= reset_n,
                              apb_request  <= gpio_apb_request,
                              apb_response => gpio_apb_response,
                              gpio_input <= gpio_input,
                              gpio_output => gpio_output,
                              gpio_output_enable => gpio_output_enable,
                              gpio_input_event => gpio_input_event
            );
        apb_target_uart_minimal uart( clk <- clk,
                                      reset_n <= reset_n,
                                      apb_request  <= uart_apb_request,
                                      apb_response => uart_apb_response,
                                      uart_rx <= uart_rx,
                                      uart_tx => uart_tx,
                                      status => uart_status
            );

        apb_target_i2c_master i2c( clk <- clk,
                                       reset_n <= reset_n,
                                       apb_request  <= i2c_apb_request,
                                       apb_response => i2c_apb_response,
                                       i2c_in  <= subsys_inputs.i2c,
                                       i2c_out => i2c_master );

        apb_target_axi4s apb_axi4s( clk <- clk,
                                    reset_n <= reset_n,
                                    apb_request  <= axi4s_apb_request,
                                    apb_response => axi4s_apb_response,
                                    tx_sram_access_req  => tx_sram_access_req,
                                    tx_sram_access_resp <= tx_sram_access_resp,
                                    rx_sram_access_req  => rx_sram_access_req,
                                    rx_sram_access_resp <= rx_sram_access_resp,
                                    rx_axi4s        <= rx_axi4s,
                                    rx_axi4s_tready => rx_axi4s_tready,
                                    tx_axi4s         => tx_axi4s,
                                    tx_axi4s_tready  <= tx_axi4s_tready );

        apb_target_analyzer apb_analyzer( apb_clock <- clk,
                                          reset_n <= reset_n,
                                          apb_request  <= anal_apb_request,
                                          apb_response => anal_apb_response,
                                          analyzer_mux_control => analyzer_mux_control,

                                          analyzer_clock <- clk,
                                          internal_signal_in <= analyzer_trace,
                             
                                          // trace_ready,
                                          // trace_done,
                                          ext_trigger_reset <= 0,
                                          ext_trigger_enable <= 0,

                                          async_trace_read_clock <- clk, // unused interface for now
                                          async_trace_read_enable <= 0
                                          // async_trace_valid_out,
                                          // async_trace_out
            );

        csr_master_apb master( clk <- clk,
                               reset_n <= reset_n,
                               apb_request <= csr_apb_request,
                               apb_response => csr_apb_response,
                               csr_request => csr_request,
                               csr_response <= csr_response_r );

    }

    /*b Dprintf/framebuffer */
    net bit dprintf_uart_txd;
    dprintf_framebuffer_instances: {
        fifo_dprintf_req_fb    = fifo_dprintf_req;
        fifo_dprintf_req_uart  = fifo_dprintf_req;
        fifo_dprintf_ack       = fifo_dprintf_ack_fb;

        if (debug.uart_src_dprintf) {
            fifo_dprintf_ack       = fifo_dprintf_ack_uart;
            fifo_dprintf_req_fb.valid  = 0;
        } else {
            fifo_dprintf_ack       = fifo_dprintf_ack_fb;
            fifo_dprintf_req_uart.valid  = 0;
        }
        apb_target_dprintf_uart apb_dprintf_uart( clk <- clk,
                                              reset_n <= reset_n,
                                              apb_request  <= dprintf_uart_apb_request,
                                              apb_response => dprintf_uart_apb_response,
                                              dprintf_req <= fifo_dprintf_req_uart,
                                              dprintf_ack => fifo_dprintf_ack_uart,
                                              uart_txd => dprintf_uart_txd );

        dprintf dprintf( clk <- clk,
                         reset_n <= reset_n,
                         dprintf_req <= fifo_dprintf_req_fb,
                         dprintf_ack => fifo_dprintf_ack_fb,
                         byte_blocked <= 0,
                         dprintf_byte => dprintf_byte
            );

        tt_display_sram_access_req = {*=0,
                                      valid = dprintf_byte.valid,
                                      address = bundle(16b0, dprintf_byte.address),
                                      write_data = bundle(56b0, dprintf_byte.data) };

        fb_sram_access_resp = {*=0};
        fb_sram_access_resp.ack   = fb_sram_access_req.valid;
        fb_sram_access_resp.valid = fb_sram_access_req.valid;
        fb_sram_access_resp.id    = fb_sram_access_req.id;

        framebuffer_teletext ftb_debug( csr_clk <- clk,
                                        sram_clk <- clk,
                                        video_clk <- video_clk,
                                        reset_n <= reset_n,
                                        video_bus => debug_video_bus,
                                        display_sram_write <= tt_display_sram_access_req,
                                        csr_select_in <= 16h2, // uses 2 selects
                                        csr_request <= csr_request,
                                        csr_response => tt_debug_framebuffer_csr_response
            );

        framebuffer_teletext ftb_vga( csr_clk <- clk,
                                      sram_clk <- clk,
                                      video_clk <- video_clk,
                                      reset_n <= reset_n,
                                      video_bus => vga_video_bus,
                                      display_sram_write <= fb_sram_access_req,
                                      csr_select_in <= 16h4, // uses 2 selects
                                      csr_request <= csr_request,
                                      csr_response => tt_vga_framebuffer_csr_response
            );

        csr_target_timeout csr_timeout(clk <- clk,
                                       reset_n <= reset_n,
                                       csr_request <= csr_request,
                                       csr_response => timeout_csr_response,
                                       csr_timeout <= 16h100 );

        csr_response  = tt_vga_framebuffer_csr_response;
        csr_response |= tt_debug_framebuffer_csr_response;
        csr_response |= timeout_csr_response;
        csr_response |= master_csr_response;
        master_csr_request = csr_request;
        csr_response_r <= csr_response;

        video_bus = vga_video_bus;
        if (debug.video_src_debug) {
            video_bus = debug_video_bus;
        }
    }

    /*b Ethernet */
    ethernet : {
        se_sram_srw_16384x32_we8 rx_mem(sram_clock <- clk,
                                     select         <= rx_sram_access_req.valid && rx_sram_access_resp.ack,
                                     read_not_write <= rx_sram_access_req.read_not_write,
                                     write_enable   <= rx_sram_access_req.byte_enable[4;0],
                                     address        <= rx_sram_access_req.address[14;0],
                                     write_data     <= rx_sram_access_req.write_data[32;0],
                                     data_out       => rx_sram_read_data );
        rx_sram_access_resp <= {*=0};
        rx_sram_access_resp.ack   <= 1;
        rx_current_sram_access.valid <= 0;
        if (rx_sram_access_req.valid && rx_sram_access_resp.ack) {
            rx_current_sram_access <= rx_sram_access_req;
        }
        if (rx_current_sram_access.valid) {
            rx_sram_access_resp.valid       <= rx_current_sram_access.read_not_write;
            rx_sram_access_resp.id          <= rx_current_sram_access.id;
            rx_sram_access_resp.data[32;0]  <= rx_sram_read_data;
        }

        se_sram_srw_16384x32_we8 tx_mem(sram_clock <- clk,
                                     select         <= tx_sram_access_req.valid && tx_sram_access_resp.ack,
                                     read_not_write <= tx_sram_access_req.read_not_write,
                                     write_enable   <= tx_sram_access_req.byte_enable[4;0],
                                     address        <= tx_sram_access_req.address[14;0],
                                     write_data     <= tx_sram_access_req.write_data[32;0],
                                     data_out       => tx_sram_read_data );
        tx_sram_access_resp <= {*=0};
        tx_sram_access_resp.ack   <= 1;
        tx_current_sram_access.valid <= 0;
        if (tx_sram_access_req.valid && tx_sram_access_resp.ack) {
            tx_current_sram_access <= tx_sram_access_req;
        }
        if (tx_current_sram_access.valid) {
            tx_sram_access_resp.valid       <= tx_current_sram_access.read_not_write;
            tx_sram_access_resp.id          <= tx_current_sram_access.id;
            tx_sram_access_resp.data[32;0]  <= tx_sram_read_data;
        }
    }
    
    /*b Subsystem outputs */
    subsystem_output_logic : {
        timer_control <= rv_timer_control;
        
        uart_rx = {*=0};
        uart_rx.rxd = subsys_inputs.uart_rx.rxd;
        if (debug.uart_src_dprintf) {
            subsys_outputs.uart_tx.txd = dprintf_uart_txd;
            subsys_outputs.uart_tx.cts = 0;
        } else {
            subsys_outputs.uart_tx= uart_tx;
        }
        subsys_outputs.reset_request = 0;
        subsys_outputs.i2c = {*=1};
        subsys_outputs.gpio_output        = gpio_output[8;8];
        subsys_outputs.gpio_output_enable = gpio_output_enable[8;8];
        gpio_input      <= 0;
        gpio_input[0]   <= subsys_inputs.i2c.scl;
        gpio_input[1]   <= subsys_inputs.i2c.sda;
        gpio_input[8;8] <= subsys_inputs.gpio_input;

        if (gpio_output_enable[0] && !gpio_output[0]) {subsys_outputs.i2c.scl = 0;}
        if (gpio_output_enable[1] && !gpio_output[1]) {subsys_outputs.i2c.sda = 0;}
        if (!i2c_master.scl) {subsys_outputs.i2c.scl = 0;}
        if (!i2c_master.sda) {subsys_outputs.i2c.sda = 0;}
    }
}
