/** Copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *   http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * @file  tb_hysteresis_switch.cdl
 * @brief Testbench for hysteresis switch
 *
 * This is a simple testbench for the hysteresis switch 
 */
/*a Includes */
include "input/hysteresis.h"

/*a External modules */
extern module se_test_harness( clock clk,
                               output bit clk_enable "Assert to enable the internal clock; this permits I/O switches to easily use a slower clock",
                               output bit input_value,
                               input bit output_value,
                               output bit[16] filter_period "Period over which to filter the input - the larger the value, the longer it takes to switch, but the more glitches are removed",
                               output bit[16] filter_level  "Value to exceed to switch output levels - the larger the value, the larger the hysteresis; must be less than filter_period"
    )
{
    timing from rising clock clk clk_enable;
    timing from rising clock clk input_value, filter_period, filter_level;
    timing to   rising clock clk output_value;
}

/*a Module */
module tb_hysteresis_switch( clock clk,
                    input bit reset_n
)
{

    /*b Nets */
    net bit clk_enable;
    net bit input_value;
    net bit output_value;
    net bit[16] filter_period;
    net bit[16] filter_level;

    /*b Instantiations */
    instantiations: {
        se_test_harness th( clk <- clk,
                            clk_enable => clk_enable,
                            input_value => input_value,
                            output_value <= output_value,
                            filter_period => filter_period,
                            filter_level => filter_level );

        hysteresis_switch hs( clk <- clk,
                              reset_n <= reset_n,
                              clk_enable <= clk_enable,
                              input_value <= input_value,
                              output_value => output_value,
                              filter_period <= filter_period,
                              filter_level <= filter_level );
    }

    /*b All done */
}
