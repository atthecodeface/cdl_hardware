/** @copyright (C) 2016-2018,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   apb_target_rv_timer.cdl
 * @brief  RISC-V compatible timer target for an APB bus
 *
 * CDL implementation of a RISC-V timer target on an APB bus,
 * supporting fractional clocks, derived from the original GIP baud
 * rate generator.
 *
 */
/*a Includes
 */
include "types/apb.h"
include "types/timer.h"
include "clocking/clock_timer_modules.h"

/*a Types */
/*t t_apb_address
 *
 * APB address map, used to decode paddr
 *
 */
typedef enum [4] {
    apb_address_timer_lower       = 0  "Bottom 32 bits of timer value; writable unless control.block_writes is high",
    apb_address_timer_upper       = 1  "Top 32 bits of timer value; writable unless control.block_writes is high",
    apb_address_comparator_lower  = 2  "Bottom 32 bits of comparator value",
    apb_address_comparator_upper  = 3  "Top 32 bits of comparator value",
} t_apb_address;

/*t t_access
 *
 * APB access that is in progress; a decode of psel and paddr
 *
 */
typedef enum [4] {
    access_none                      "No access being performed",
    access_write_timer_lower         "Write to bottom 32 bits of timer",
    access_write_timer_upper         "Write to top 32 bits of timer",
    access_read_timer_lower          "Read of bottom 32 bits of timer",
    access_read_timer_upper          "Read of top 32 bits of timer",
    access_write_comparator_lower    "Write to bottom 32 bits of comparator",
    access_write_comparator_upper    "Write to top 32 bits of comparator",
    access_read_comparator_lower     "Read of bottom 32 bits of comparator",
    access_read_comparator_upper     "Read of top 32 bits of comparator"
} t_access;

/*t t_timer_combs
 *
 */
typedef struct {
    bit[33] lower_t_minus_c  "Difference between timer and comparator lower halves, with borrow bit";
    bit[33] upper_t_minus_c  "Difference between timer and comparator upper halves, with borrow bit";
    t_timer_control timer_control "Timer control including write ability";
} t_timer_combs;

/*t t_timer_state
 *
 */
typedef struct {
    bit[32] comparator_lower       "Lower 32-bits of comparator value";
    bit[32] comparator_upper       "Upper 32-bits of comparator value";
    bit     upper_eq               "Asserted if comparator_upper==timer_upper; pipelined by 1 cycle";
    bit     upper_ge               "Asserted if comparator_upper>=timer_upper; pipelined by 1 cycle";
    bit     lower_eq               "Asserted if comparator_lower==timer_lower; pipelined by 1 cycle";
    bit     lower_ge               "Asserted if comparator_lower>=timer_lower; pipelined by 1 cycle";
    bit     comparator_exceeded    "Asserted if comparator>timer; pipelined by 2 cycles";
} t_timer_state;

/*a Module */
module apb_target_rv_timer( clock clk             "System clock",
                            input bit reset_n     "Active low reset",
                            input t_timer_control timer_control "Control of the timer", 

                            input  t_apb_request  apb_request  "APB request",
                            output t_apb_response apb_response "APB response",

                            output t_timer_value  timer_value
    )
"""
RISC-V compatible timer with an APB interface.

This is a monotonically increasing 64-bit timer with a 64-bit comparator.

"""
{
    /*b Clock and reset */
    default clock clk;
    default reset active_low reset_n;

    /*b Decode APB interface */
    clocked t_access access=access_none   "Access being performed by APB";

    /*b Timer state */
    clocked t_timer_state timer_state= {*=0} "State of the timer and comparator";
    comb    t_timer_combs timer_combs        "Combinatorial decode of timer state and controls";

    /*b APB interface */
    apb_interface_logic """
    The APB interface is decoded to @a access when @p psel is asserted
    and @p penable is deasserted - this is the first cycle of an APB
    access. This permits the access type to be registered, so that the
    APB @p prdata can be driven from registers, and so that writes
    will occur correctly when @p penable is asserted.

    The APB read data @p prdata can then be generated based on @a
    access.
    """ : {
        /*b Decode access */
        access <= access_none;
        part_switch (apb_request.paddr[4;0]) {
        case apb_address_timer_lower: {
            access <= (apb_request.pwrite && !timer_control.block_writes) ? access_write_timer_lower : access_read_timer_lower;
        }
        case apb_address_timer_upper: {
            access <= (apb_request.pwrite && !timer_control.block_writes) ? access_write_timer_upper : access_read_timer_upper;
        }
        case apb_address_comparator_lower: {
            access <= apb_request.pwrite ? access_write_comparator_lower : access_read_comparator_lower;
        }
        case apb_address_comparator_upper: {
            access <= apb_request.pwrite ? access_write_comparator_upper : access_read_comparator_upper;
        }
        }
        if (!apb_request.psel || apb_request.penable) {
            access <= access_none;
        }

        /*b Handle APB read data */
        apb_response = {*=0, pready=1};
        part_switch (access) {
        case access_read_timer_lower: {
            apb_response.prdata = timer_value_without_irq.value[32; 0];
        }
        case access_read_timer_upper: {
            apb_response.prdata = timer_value_without_irq.value[32;32];
        }
        case access_read_comparator_lower: {
            apb_response.prdata = timer_state.comparator_lower;
        }
        case access_read_comparator_upper: {
            apb_response.prdata = timer_state.comparator_upper;
        }
        }

        /*b All done */
    }

    /*b Handle the timer and comparator */
    net t_timer_value  timer_value_without_irq;
    timer_logic """
    The @a timer value can be reset or it may count on a tick, or it
    may just hold its value. Furthermore, it may be writable (the
    RISC-V spec seems to require this, but it defeats the purpose of a
    global clock if there are many of these in a system that are not
    at the same global value).

    The comparison logic operates over two clock ticks. In the first
    clock tick the upper and lower halves are subtracted to provide
    'greater-or-equal' comparisons and 'equality' comparison; these
    bits are recorded, and in a second clock tick they are combined
    and a result is generated and registered.
    """: {
        /*b Comparison logic */
        timer_combs.lower_t_minus_c = bundle(1b0, timer_value_without_irq.value[32; 0]) - bundle(1b0, timer_state.comparator_lower);
        timer_combs.upper_t_minus_c = bundle(1b0, timer_value_without_irq.value[32;32]) - bundle(1b0, timer_state.comparator_upper);
        timer_state.upper_ge <= (!timer_combs.upper_t_minus_c[32]);
        timer_state.upper_eq <= (timer_combs.upper_t_minus_c==0);
        timer_state.lower_ge <= (!timer_combs.lower_t_minus_c[32]);
        timer_state.lower_eq <= (timer_combs.lower_t_minus_c==0);
        timer_state.comparator_exceeded <= 0;
        if (timer_state.upper_eq) {
            timer_state.comparator_exceeded <= timer_state.lower_ge && !timer_state.lower_eq;
        } elsif (timer_state.upper_ge) {
            timer_state.comparator_exceeded <= 1;
        }

        /*b Write to timer value */
        timer_combs.timer_control = timer_control;
        if (access==access_write_timer_lower) {
            timer_combs.timer_control.synchronize[0] = 1;
            timer_combs.timer_control.synchronize_value[32;0] = apb_request.pwdata;
        }
        if (access==access_write_timer_upper) {
            timer_combs.timer_control.synchronize[1] = 1;
            timer_combs.timer_control.synchronize_value[32;32] = apb_request.pwdata;
        }

        /*b Instantiate the timer */
        clock_timer timer(clk <- clk,
                          reset_n <= reset_n,
                          timer_control <= timer_combs.timer_control,
                          timer_value   => timer_value_without_irq );
        
        /*b Write to comparator and timer value */
        if (access==access_write_comparator_lower) {
            timer_state.comparator_lower <= apb_request.pwdata;
        }
        if (access==access_write_comparator_upper) {
            timer_state.comparator_upper <= apb_request.pwdata;
        }

        /*b Drive outputs */
        timer_value      = timer_value_without_irq;
        timer_value.irq  = timer_state.comparator_exceeded;
    }

    /*b Done
     */
}

/*a Editor preferences and notes
mode: c ***
c-basic-offset: 4 ***
c-default-style: (quote ((c-mode . "k&r") (c++-mode . "k&r"))) ***
outline-regexp: "/\\\*a\\\|[\t ]*\/\\\*[b-z][\t ]" ***
*/
