/** Copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *   http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * @file  teletext.cdl
 * @brief CDL implementation of a teletext decoder
 *
 * This is an implementaion of the core of a teletext decoder, for
 * arbitrary sized teletext output displays.
 *
 * The output is supplied at 12 pixels per clock (one character width)
 * The input is a byte of per clock of character data.
 *
 * The implementation does not currently support double width or
 * double height characters.
 *
 */
/*a Includes */
include "teletext.h"

/*a Types */
typedef bit[3] t_color;
/*t t_character_state */
typedef struct {
    bit[3] background_color;
    bit[3] foreground_color;
    bit    held_character;
    bit    flashing;
    bit    text_mode;
    bit    contiguous_graphics;
    bit    dbl_height;
    bit    hold_graphics;
    bit    reset_held_graphics;
} t_character_state;

/*t t_load_state */
typedef struct {
    t_teletext_character character;
} t_load_state;
constant integer flashing_on_count=10;
constant integer max_flashing_count=40;

/*t t_timing_state */
typedef struct {
    bit[5] scanline;
    bit last_scanline;
    t_teletext_timings timings;
    bit[6] flashing_counter; // 50 fields per second, 3/4 second, max of ~40, flash on at 10
    bit    flash_on;
    bit    scanline_displayed "Asserted if there has been a valid character in the scanline";
} t_timing_state;

/*t t_teletext_combs */
typedef struct {
    t_character_state next_character_state;
    t_character_state current_character_state;
    bit can_be_replaced_with_hold;
    bit[5] pixel_scanline;
} t_teletext_combs;

/*t t_teletext_state */
typedef struct {
    t_teletext_character character "Used for graphics decode";
    t_character_state character_state;
    bit row_contains_dbl_height;
    bit last_row_contained_dbl_height;
} t_teletext_state;

/*t t_pixel_combs */
typedef struct {
    bit[10] rom_scanline_data;
    bit[12] graphics_data;
    bit[12] smoothed_scanline_data;
    bit[5] diagonal_0;
    bit[5] diagonal_1;
    bit[5] diagonal_2;
    bit[5] diagonal_3;
} t_pixel_combs;

/*t t_output_state */
typedef struct {
    t_character_state character_state;
    bit[12] held_graphics_data;
    t_color[12] colors;
    bit valid;
} t_output_state;

/*a Module teletext */
module teletext( clock clk     "Character clock",
                 input bit reset_n,
                 input t_teletext_character    character  "Parallel character data in, with valid signal",
                 input t_teletext_timings      timings    "Timings for the scanline, row, etc",
                 output t_teletext_rom_access  rom_access "Teletext ROM access",
                 input bit[45]                 rom_data   "Teletext ROM data, valid in cycle after rom_access",
                 output t_teletext_pixels pixels       "Output pixels, two clock ticks delayed from clk in"
       )
    /*b Documentation */
"""
Teletext characters are displayed from a 12x20 grid.
The ROM characters have two background rows, and then are displayed with 2 background pixels on the left, and then 10 pixels from the ROM
The ROM is actually 5x9, and it is doubled to 10x18
Doubling without smoothing can be achieved be true doubling

A simple smoothing can be performed for a pixel depending on its NSEW neighbors:

  |NN|
  |NN|
WW|ab|EE
WW|cd|EE
  |SS|
  |SS|

a is filled if the pixel is filled itself, or if N&W
b is filled if the pixel is filled itself, or if N&E
c is filled if the pixel is filled itself, or if S&W
d is filled if the pixel is filled itself, or if S&E

Hence one would get:
..|**|**|**|..|
..|**|**|**|..|
---------------
**|..|..|**|**|
**|..|..|**|**|
---------------
..|**|..|..|**|
..|**|..|..|**|

smoothed to:
..|**|**|**|..|
.*|**|**|**|*.|
---------------
**|*.|.*|**|**|
**|*.|..|**|**|
---------------
.*|**|..|.*|**|
..|**|..|..|**|

Or, without intervening lines:
..******..
..******..
**....****
**....****
..**....**
..**....**

smoothed to:
..******..
.********.
***..*****
***...****
.***...***
..**....**

So for even scanlines ('a' and 'b') the smoother needs row n and row n-1.
a is set if n[x] or n[x-left]&(n-1)[x]
b is set if n[x] or n[x-right]&(n-1)[x]

For odd scanlines ('c' and 'd') the smoother needs row n and row n+1.
c is set if n[x] or n[x-left]&(n+1)[x]
d is set if n[x] or n[x-right]&(n+1)[x]

This method has the unfortunate impact of smoothing two crossing lines, such as a plus:
....**....     ....**....
....**....     ....**....
....**....     ....**....
....**....     ...****...
**********     **********
**********     **********
....**....     ...****...
....**....     ....**....
....**....     ....**....
....**....     ....**....

Hence a better smoothing can be performed for a pixel depending on all its neighbors:

NW|NN|NE
  |NN|
WW|ab|EE
WW|cd|EE
  |SS|
SW|SS|SE

a is filled if the pixel is filled itself, or if (N&W) but not NW
b is filled if the pixel is filled itself, or if (N&E) but not NE
c is filled if the pixel is filled itself, or if (S&W) but not SW
d is filled if the pixel is filled itself, or if (S&E) but not SE

Hence one would get:
..|**|**|**|..|
..|**|**|**|..|
---------------
**|..|..|**|**|
**|..|..|**|**|
---------------
..|**|..|..|**|
..|**|..|..|**|

smoothed to:
..|**|**|**|..|
.*|**|**|**|..|
---------------
**|*.|..|**|**|
**|*.|..|**|**|
---------------
.*|**|..|..|**|
..|**|..|..|**|

Or, without intervening lines:
..******..
..******..
**....****
**....****
..**....**
..**....**

smoothed to:
..******..
.*******..
***...****
***...****
.***....**
..**....**

So for even scanlines ('a' and 'b') the smoother needs row n and row n-1.
a is set if n[x] or (n[x-left]&(n-1)[x]) &~ (n-1)[x-left]
b is set if n[x] or (n[x-right]&(n-1)[x]) &~ (n-1)[x-right]

For odd scanlines ('c' and 'd') the smoother needs row n and row n+1.
c is set if n[x] or (n[x-left]&(n+1)[x]) &~ (n+1)[x-left]
d is set if n[x] or (n[x-right]&(n+1)[x]) &~ (n+1)[x-left]

Graphics characters are 6 blobs on a 6x10 grid (contiguous, separated):
000111 .00.11
000111 .00.11
000111 ......
222333 .22.33
222333 .22.33
222333 .22.33
222333 ......
444555 .44.55
444555 .44.55
444555 ......

"""
{
    /*b Defaults */
    default reset active_low reset_n;
    default clock clk;
    clocked t_load_state      load_state = {*=0};
    clocked t_timing_state    timing_state = {*=0};
    clocked t_teletext_state  teletext_state = {*=0};
    clocked t_teletext_rom_access  rom_access = {*=0};
    comb    t_teletext_combs  teletext_combs;
    comb    t_pixel_combs     pixel_combs;
    clocked t_output_state output_state={*=0};

    /*b Timing control and load_state stage */
    scanline_and_loading """
    """: {
        load_state.character <= character;

        rom_access.select <= 0;
        if (character.valid) {
            rom_access <= {select=1,
                    address = character.character};
        }

        timing_state.timings <= timings;
        timing_state.scanline <= timing_state.scanline+2;
        if (timing_state.timings.interpolate_vertical == tvi_all_scanlines) {
            timing_state.scanline <= timing_state.scanline+1;
        }
        if (timing_state.last_scanline || timings.first_scanline_of_row) {
            timing_state.scanline <= 0;
            if (timing_state.timings.interpolate_vertical == tvi_odd_scanlines) {
                timing_state.scanline <= 1;
            }
        }
        timing_state.last_scanline <= 0;
        if (timing_state.scanline==19) {
            timing_state.last_scanline <= 1;
        }
        if ((timing_state.scanline==18) && (timing_state.timings.interpolate_vertical == tvi_even_scanlines)){
            timing_state.last_scanline <= 1;
        }

        if (!timings.first_scanline_of_row && !timings.end_of_scanline) {
            timing_state.scanline <= timing_state.scanline;
        }
        if (!timing_state.scanline_displayed) {
            timing_state.scanline <= timing_state.scanline;
        }
        if (timings.end_of_scanline) {
            timing_state.scanline_displayed <= 0;
        }
        if (load_state.character.valid) {
            timing_state.scanline_displayed <= 1;
        }

        if (timings.restart_frame) {
            timing_state.flashing_counter <= timing_state.flashing_counter+1;
            if (timing_state.flashing_counter==flashing_on_count) {
                timing_state.flash_on <= 1;
            }
            if (timing_state.flashing_counter==max_flashing_count) {
                timing_state.flashing_counter <= 0;
                timing_state.flash_on <= 0;
            }
        }
    }

    /*b Teletext control decode */
    teletext_control_decode """
    Decode the 'load_state' character if a control character; handle the state of the line (colors, graphics, etc)
    """: {
        /*b Decode current character while reading its contents from ROM
          note that steady, normal size, conceal, contiguous, separated, black background, new background, hold are 'set-at'
          rest are 'set-after'.
          'set-at' means it takes immediate effect for this character, 'set-after' just for the following characters
         */
        teletext_combs.next_character_state    = teletext_state.character_state;
        teletext_combs.current_character_state = teletext_state.character_state;
        teletext_combs.can_be_replaced_with_hold = 1;
        teletext_combs.current_character_state.reset_held_graphics = 0;
        part_switch (load_state.character.character) {
        case 0: { // probably also the other un-interpreted <32 characters...
            teletext_combs.can_be_replaced_with_hold = 1;
        }
        case 1,2,3,4,5,6,7: {
            teletext_combs.next_character_state.foreground_color = load_state.character.character[3;0];
            teletext_combs.next_character_state.text_mode = 1;
            teletext_combs.current_character_state.hold_graphics = 0; // Note that this is leaving mosaics mode
            teletext_combs.next_character_state.hold_graphics = 0; // immediately... hence no hold for this
            teletext_combs.current_character_state.reset_held_graphics = !teletext_state.character_state.text_mode;
        }
        case 8: { teletext_combs.next_character_state.flashing = 1; }
        case 9: { // steady is set-at
            teletext_combs.current_character_state.flashing = 0;
            teletext_combs.next_character_state.flashing = 0;
            // does this reset the held graphics?
        }
        case 17,18,19,20,21,22,23: {
            teletext_combs.next_character_state.foreground_color = load_state.character.character[3;0];
            teletext_combs.next_character_state.text_mode = 0;
            teletext_combs.current_character_state.reset_held_graphics = teletext_state.character_state.text_mode;
            // does this reset the held graphics?
        }
        case 12: { // normal size is set-at
            teletext_combs.current_character_state.dbl_height = 0;
            teletext_combs.next_character_state.dbl_height    = 0;
            teletext_combs.current_character_state.reset_held_graphics = 1;
            // does this reset the held graphics?
        }
        case 13: { // double height is set-after
            teletext_combs.current_character_state.reset_held_graphics = 1;
            teletext_combs.next_character_state.dbl_height = 1;
            // does this reset the held graphics?
        }
        case 25: { // contiguous graphics is set-at
            teletext_combs.current_character_state.contiguous_graphics = 1;
            teletext_combs.next_character_state.contiguous_graphics = 1;
        }
        case 26: { // separated graphics is set-at
            teletext_combs.current_character_state.contiguous_graphics = 0;
            teletext_combs.next_character_state.contiguous_graphics = 0;
        }
        case 28: { // black background is set-at
            teletext_combs.current_character_state.background_color = 0;
            teletext_combs.next_character_state.background_color = 0;
        }
        case 29: { // new background is set-at
            teletext_combs.current_character_state.background_color = teletext_state.character_state.foreground_color;
            teletext_combs.next_character_state.background_color    = teletext_state.character_state.foreground_color;
        }
        case 30: { // hold mode is set-at
            teletext_combs.current_character_state.hold_graphics = 1; // note that a held character is the last graphics character INCLUDING separated or not
            teletext_combs.next_character_state.hold_graphics = 1;
        }
        case 31: { // release graphics is set-after
            teletext_combs.next_character_state.hold_graphics = 0;
        }
        default: {
            teletext_combs.can_be_replaced_with_hold = 0;
        }
        }

        /*b Determine scanline - using double height if necessary */
        teletext_combs.pixel_scanline = timing_state.scanline;
        if (teletext_state.character_state.dbl_height) {
            teletext_combs.pixel_scanline = bundle(1b0,timing_state.scanline[4;1]);
            if (teletext_state.last_row_contained_dbl_height) {
                teletext_combs.pixel_scanline = teletext_combs.pixel_scanline + 10;
            }
        }

        /*b Handle change of control state at end of character */
        teletext_state.character.valid <= 0;
        if (load_state.character.valid) {
            teletext_state.character <= load_state.character;
            teletext_state.character_state  <= teletext_combs.next_character_state;
            if (teletext_combs.current_character_state.dbl_height) {
                teletext_state.row_contains_dbl_height <= 1;
            }
        }

        /*b Handle reset of control state at end of scanline */
        if (timing_state.timings.end_of_scanline) {
            teletext_state.character_state.background_color <= 0;
            teletext_state.character_state.foreground_color <= 3b111;
            teletext_state.character_state.held_character <= 0;
            teletext_state.character_state.flashing <= 0;
            teletext_state.character_state.dbl_height <= 0;
            teletext_state.character_state.text_mode <= 1;
            teletext_state.character_state.hold_graphics <= 0;
            teletext_state.character_state.contiguous_graphics <= 1;
        }

        /*b Handle reset of control state at end of character row */
        if (timing_state.timings.end_of_scanline && timing_state.last_scanline) {
            teletext_state.last_row_contained_dbl_height <= teletext_state.row_contains_dbl_height ^ teletext_state.last_row_contained_dbl_height;
            teletext_state.row_contains_dbl_height <= 0;
        }

        /*b Handle reset of control state at end of field */
        if (timing_state.timings.restart_frame) {
            teletext_state.last_row_contained_dbl_height <= 0;
            teletext_state.row_contains_dbl_height <= 0;
        }
    }

    /*b Character ROM fetch and pixel data generation - in same stage as control decode */
    character_rom_and_pixel_generation """
    """: {
        /*b Select scanline of ROM data for pixel */
        full_switch (teletext_combs.pixel_scanline[4;1]) { //scanline_of_character changes every scanline, so no need to have a pixel pipeline stage version
        case 0: { pixel_combs.rom_scanline_data = bundle(rom_data[5;0],5b0); }
        case 1: { pixel_combs.rom_scanline_data = rom_data[10;0]; }
        case 2: { pixel_combs.rom_scanline_data = rom_data[10;5]; }
        case 3: { pixel_combs.rom_scanline_data = rom_data[10;10]; }
        case 4: { pixel_combs.rom_scanline_data = rom_data[10;15]; }
        case 5: { pixel_combs.rom_scanline_data = rom_data[10;20]; }
        case 6: { pixel_combs.rom_scanline_data = rom_data[10;25]; }
        case 7: { pixel_combs.rom_scanline_data = rom_data[10;30]; }
        case 8: { pixel_combs.rom_scanline_data = rom_data[10;35]; }
        default: { pixel_combs.rom_scanline_data = bundle(5b0,rom_data[5;40]); } // 9, and catch-all
        }

        /*b Smoothe ROM data for pixel */
        pixel_combs.diagonal_0 = pixel_combs.rom_scanline_data[5;5] & bundle(pixel_combs.rom_scanline_data[4;0], 1b0);
        pixel_combs.diagonal_1 = pixel_combs.rom_scanline_data[5;5] & bundle(1b0,pixel_combs.rom_scanline_data[4;1]);
        pixel_combs.diagonal_2 = pixel_combs.rom_scanline_data[5;0] & bundle(pixel_combs.rom_scanline_data[4;5], 1b0);
        pixel_combs.diagonal_3 = pixel_combs.rom_scanline_data[5;0] & bundle(1b0,pixel_combs.rom_scanline_data[4;6]);

        pixel_combs.diagonal_0 = pixel_combs.diagonal_0 &~ bundle(pixel_combs.rom_scanline_data[4;5], 1b0);
        pixel_combs.diagonal_1 = pixel_combs.diagonal_1 &~ bundle(1b0,pixel_combs.rom_scanline_data[4;6]);
        pixel_combs.diagonal_2 = pixel_combs.diagonal_2 &~ bundle(pixel_combs.rom_scanline_data[4;0], 1b0);
        pixel_combs.diagonal_3 = pixel_combs.diagonal_3 &~ bundle(1b0,pixel_combs.rom_scanline_data[4;1]);
        if (!teletext_combs.pixel_scanline[0]) {
            pixel_combs.smoothed_scanline_data = bundle( 2b0,
                                                         pixel_combs.rom_scanline_data[4]|pixel_combs.diagonal_1[4],
                                                         pixel_combs.rom_scanline_data[4]|pixel_combs.diagonal_0[4],
                                                         pixel_combs.rom_scanline_data[3]|pixel_combs.diagonal_1[3],
                                                         pixel_combs.rom_scanline_data[3]|pixel_combs.diagonal_0[3],
                                                         pixel_combs.rom_scanline_data[2]|pixel_combs.diagonal_1[2],
                                                         pixel_combs.rom_scanline_data[2]|pixel_combs.diagonal_0[2],
                                                         pixel_combs.rom_scanline_data[1]|pixel_combs.diagonal_1[1],
                                                         pixel_combs.rom_scanline_data[1]|pixel_combs.diagonal_0[1],
                                                         pixel_combs.rom_scanline_data[0]|pixel_combs.diagonal_1[0],
                                                         pixel_combs.rom_scanline_data[0]|pixel_combs.diagonal_0[0]
                );
        } else {
            pixel_combs.smoothed_scanline_data = bundle( 2b0,
                                                         pixel_combs.rom_scanline_data[9]|pixel_combs.diagonal_3[4],
                                                         pixel_combs.rom_scanline_data[9]|pixel_combs.diagonal_2[4],
                                                         pixel_combs.rom_scanline_data[8]|pixel_combs.diagonal_3[3],
                                                         pixel_combs.rom_scanline_data[8]|pixel_combs.diagonal_2[3],
                                                         pixel_combs.rom_scanline_data[7]|pixel_combs.diagonal_3[2],
                                                         pixel_combs.rom_scanline_data[7]|pixel_combs.diagonal_2[2],
                                                         pixel_combs.rom_scanline_data[6]|pixel_combs.diagonal_3[1],
                                                         pixel_combs.rom_scanline_data[6]|pixel_combs.diagonal_2[1],
                                                         pixel_combs.rom_scanline_data[5]|pixel_combs.diagonal_3[0],
                                                         pixel_combs.rom_scanline_data[5]|pixel_combs.diagonal_2[0]
                );
        }
        if (!timing_state.timings.smoothe) {
            pixel_combs.smoothed_scanline_data = bundle( 2b0,
                                                         pixel_combs.rom_scanline_data[4],pixel_combs.rom_scanline_data[4],
                                                         pixel_combs.rom_scanline_data[3],pixel_combs.rom_scanline_data[3],
                                                         pixel_combs.rom_scanline_data[2],pixel_combs.rom_scanline_data[2],
                                                         pixel_combs.rom_scanline_data[1],pixel_combs.rom_scanline_data[1],
                                                         pixel_combs.rom_scanline_data[0],pixel_combs.rom_scanline_data[0] );
        }

        /*b Generate graphcis data */
        pixel_combs.graphics_data = 12h00;
        full_switch (teletext_combs.pixel_scanline[4;1]) {
        case 0, 1, 2: {
            pixel_combs.graphics_data = (teletext_state.character.character[0]?12hfc0:12h0) | (teletext_state.character.character[1]?12h03f:12h0);
        }
        case 7,8,9: {
            pixel_combs.graphics_data = (teletext_state.character.character[4]?12hfc0:12h0) | (teletext_state.character.character[6]?12h03f:12h0);
        }
        default: {
            pixel_combs.graphics_data = (teletext_state.character.character[2]?12hfc0:12h0) | (teletext_state.character.character[3]?12h03f:12h0);
        }
        }
        if (!output_state.character_state.contiguous_graphics) {
            pixel_combs.graphics_data[2;10] = 2b00;
            pixel_combs.graphics_data[2; 4]  = 2b00;
            part_switch (teletext_combs.pixel_scanline[4;1]) {
            case 2, 6, 9: {pixel_combs.graphics_data = 0;}
            }
        }

        /*b Override character ROM if in graphics mode or held*/
        if (!output_state.character_state.text_mode) {
            if (teletext_state.character.character[5]) {
                pixel_combs.smoothed_scanline_data = pixel_combs.graphics_data;
                output_state.held_graphics_data <= pixel_combs.graphics_data;
            }
        }
        if (output_state.character_state.hold_graphics && (teletext_state.character.character[2;5]==0)) {
            pixel_combs.smoothed_scanline_data = output_state.held_graphics_data;
        }

        if (timing_state.timings.end_of_scanline) {
            output_state.held_graphics_data <= 0;
        }
        if (output_state.character_state.reset_held_graphics) {
            output_state.held_graphics_data <= 0;
        }
    }

    /*b Character pixel generation, in pixel pipeline stage and outputs */
    character_pixel_generation """
    Get two scanlines - current and next (next of 0 if none)
    """: {
        output_state.character_state <= teletext_combs.current_character_state;
        output_state.valid <= teletext_state.character.valid;

        pixels.red = 0;
        pixels.blue = 0;
        pixels.green = 0;
        for (i; 12) {
            output_state.colors[i] <= pixel_combs.smoothed_scanline_data[i] ? output_state.character_state.foreground_color : output_state.character_state.background_color;
        }
        for (i; 12) {
            pixels.red[i]   = output_state.colors[i][0];
            pixels.green[i] = output_state.colors[i][1];
            pixels.blue[i]  = output_state.colors[i][2];
        }
        pixels.valid = output_state.valid;
        pixels.last_scanline = timing_state.last_scanline;
    }

    /*b All done */
}
