/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   async_reduce.cdl
 * @brief  Reduce a bus from one clock domain to another
 *
 */
/*a Includes */
include "technology/sync_modules.h"

/*a Constants */
constant integer input_width  = 4;
constant integer double_sr    = 0;
constant integer output_width = 60;
constant integer shift_register_width = (double_sr+1)*output_width;
constant integer shift_right = 1;
constant integer cycles = shift_register_width / input_width;
constant integer counter_size = sizeof(cycles);

/*a Types */
/*t t_sr */
typedef bit[shift_register_width] t_sr;

/*t t_data_in_state */
typedef struct {
    bit[counter_size] counter;
    t_sr shift_register;
    t_sr data_out;
    bit  data_valid_toggle;
} t_data_in_state;

/*t t_data_out_state */
typedef struct {
    bit    last_valid_toggle;
    t_sr   data_out;
    bit[2] data_out_valid   "One bit for each half of the shift register - if not doubled, then always 0 or 3";
} t_data_out_state;

/*a Module
 */
module generic_async_reduce( clock clk_in "Clock associated with data_in",
                             clock clk_out "Clock associated with data_out",
                             input bit reset_n,
                             input bit valid_in,
                             input bit[input_width] data_in,
                             output bit               valid_out,
                             output bit[output_width] data_out
    )
"""
Take in a bus of @a input_width bits, and use a shift register to
shift into an output (configurable direction) of @a output_width bits
Then synchronize to the output clock domain.

If @a shift_right then the data is shifted right as it comes in - older data is at the right
Else older data is at the left

The shift register can be configured to be twice the width of the output data, with a single
synchronization used for that double width.

The synchronization between clk_in and clk_out is a tech synchronizer of a toggle.
Assuming clk_in rises at time 0 generating a toggle, the first flop of the synchronizer
occurs on clk_out at up to a whole clk_out period later; the second flop of the synchronizer
occurs up to two clk_out periods later; the data is captured on the next edge (when sync != last
toggle) - i.e. three clk_out periods later.

Hence the design works if clk_out period*3 is less than clk_in period * shift_register_width/input_width.

A shift register which is double the size of the output_width can meet this too.

This permits a 4-bit input at 312.5MHz (3.2ns period) to transfer to a 125MHz domain (8ns period)
(clk_out/clk_in periods of 2.5) with a shift register width of >30 bits.
Using a double shift register of 56 bits yields two consecutive output cycles every 14 input clocks,
or 44.8ns; hence two out of every 5.6 cycles.

"""
{
    /*b Clock in domain */
    default reset active_low reset_n;
    default clock clk_in;
    clocked t_data_in_state data_in_state={*=0};
    clk_in_domain: {
        if (shift_right) {
            data_in_state.shift_register <= data_in_state.shift_register >> input_width;
            data_in_state.shift_register[input_width;shift_register_width-input_width] <= data_in;
        } else {
            data_in_state.shift_register <= data_in_state.shift_register << input_width;
            data_in_state.shift_register[input_width;0] <= data_in;
        }
        data_in_state.counter <= data_in_state.counter-1;
        if (data_in_state.counter==0) {
            data_in_state.counter <= cycles-1;
            data_in_state.data_out <= data_in_state.shift_register;
            data_in_state.data_valid_toggle <= !data_in_state.data_valid_toggle;
        }
        if (!valid_in) {
            data_in_state <= data_in_state;
        }
    }

    /*b Clock out domain */
    default reset active_low reset_n;
    default clock clk_out;
    net bit clk_out_valid_toggle_sync;
    clocked t_data_out_state data_out_state={*=0};
    clk_out_domain: {
        tech_sync_bit clk_out_toggle_sync(clk <- clk_out,
                                           reset_n <= reset_n,
                                           d <= data_in_state.data_valid_toggle,
                                           q => clk_out_valid_toggle_sync );
        data_out_state.last_valid_toggle <= clk_out_valid_toggle_sync;
        data_out_state.data_out_valid <= 0;
        if (double_sr && data_out_state.data_out_valid[0]) {
            data_out_state.data_out_valid <= data_out_state.data_out_valid>>1;
            data_out_state.data_out       <= data_out_state.data_out>>output_width;
        }
        if (data_out_state.last_valid_toggle != clk_out_valid_toggle_sync) {
            data_out_state.data_out       <= data_in_state.data_out;
            data_out_state.data_out_valid <= 3;
            if (double_sr && !shift_right) {
                for (i; 1+double_sr) { // swap halves if double and shift left
                    data_out_state.data_out[output_width;output_width*i] <= data_in_state.data_out[output_width;(double_sr-i)*output_width];
                }
            }
        }
        valid_out = data_out_state.data_out_valid[0];
        data_out[output_width;0]  = data_out_state.data_out[output_width;0];
    }
}
