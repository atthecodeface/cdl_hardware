/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   apb_target_timer.cdl
 * @brief  Simple timer target for an APB bus
 *
 * CDL implementation of a simple timer target on an APB bus, derived
 * from an original GIP version.
 *
 */
/*a Includes
 */
include "types/apb.h"
include "boards/de1_cl/de1_cl_types.h"

/*a Types */
/*t t_apb_address
 *
 * APB address map, used to decode paddr
 */
typedef enum [5] {
    apb_address_state = 0    "Address for accessing the state of the inputs",
    apb_address_dials = 1    "Address for accessing the state of the two rotary dials",
} t_apb_address;

/*t t_access
 *
 * APB access that is in progress; a decode of psel and paddr
 */
typedef enum [3] {
    access_none,
    access_read_state,
    access_read_dials,
} t_access;

/*t t_input_state
 *
 * Clock divider and LED contents
 *
 */
typedef struct
{
    t_de1_cl_user_inputs user_inputs;
    bit    inputs_changed "Asserted if inputs have changed since last read";
    bit[8] left_dial_position;
    bit[8] right_dial_position;
} t_input_state;

/*a Module */
module apb_target_de1_cl_inputs( clock clk         "System clock",
                                 input bit reset_n "Active low reset",

                                 input  t_apb_request  apb_request  "APB request",
                                 output t_apb_response apb_response "APB response",

                                 input t_de1_cl_user_inputs    user_inputs
    )
"""
This module provides an APB target to get the status of inputs for the
Cambridge University DE1-SOC daughterboard.

The CL DE1-SOC daughterboard contains a joystick, a diamond of four
buttons, two rotary dials, and apparently a temperature alarm and
touchpanel intrerrupt (the latter two I have not used as yet).

Two registers are provided. The first is the state register,

Bits     | Meaning
---------|---------
31       | Inputs changed since last read of state
5;26     | zero
25       | temperature alarm
24       | touchpanel interrupt
6;18     | zero
17       | right rotary dial is pressed in
16       | left rotary dial is pressed in
3;13     | zero
12       | joystick is being pressed
11       | joystick is being pushed right
10       | joystick is being pushed left
9        | joystick is being pushed down
8        | joystick is being pushed up
4;4      | zero
3        | diamond y (top black button) is being pressed
2        | diamond x (left blue button) is being pressed
1        | diamond b (right red button) is being pressed
0        | diamond a (bottom green button) is being pressed

The second register relates just to the rotary dials; the hardware
keeps track of directional impulses to provide an 8-bit 'rotary value'
for each dial.

Bits     | Meaning
---------|---------
31       | Inputs changed since last read of state
13;18     | zero
17       | right rotary dial is pressed in
16       | left rotary dial is pressed in
8;8      | right rotary dial position (decremented on anticlockwise, incremented on clockwise)
8;0      | left rotary dial position (decremented on anticlockwise, incremented on clockwise)
"""
{
    /*b Clock and reset */
    default clock clk;
    default reset active_low reset_n;

    /*b Decode APB interface */
    clocked t_access access=access_none   "Access being performed by APB";

    /*b Timer state */
    clocked t_input_state input_state={*=0};

    /*b APB interface */
    apb_interface_logic """
    The APB interface is decoded to @a access when @p psel is asserted
    and @p penable is deasserted - this is the first cycle of an APB
    access. This permits the access type to be registered, so that the
    APB @p prdata can be driven from registers, and so that writes
    will occur correctly when @p penable is asserted.

    The APB read data @p prdata can then be generated based on @a
    access.
    """ : {
        /*b Decode access */
        access <= access_none;
        part_switch (apb_request.paddr[3;0]) {
        case apb_address_state: {
            access <= apb_request.pwrite ? access_none : access_read_state;
        }
        case apb_address_dials: {
            access <= apb_request.pwrite ? access_none : access_read_dials;
        }
        }
        if (!apb_request.psel || apb_request.penable) {
            access <= access_none;
        }

        /*b Handle APB read data */
        apb_response = {*=0, pready=1};
        part_switch (access) {
        case access_read_state: {
            apb_response.prdata = bundle( input_state.inputs_changed,
                                          5b0,
                                          input_state.user_inputs.temperature_alarm,
                                          input_state.user_inputs.touchpanel_irq,
                                          6b0,
                                          input_state.user_inputs.right_dial.pressed,
                                          input_state.user_inputs.left_dial.pressed,
                                          3b0,
                                          input_state.user_inputs.joystick.c,
                                          input_state.user_inputs.joystick.r,
                                          input_state.user_inputs.joystick.l,
                                          input_state.user_inputs.joystick.d,
                                          input_state.user_inputs.joystick.u,
                                          4b0,
                                          input_state.user_inputs.diamond.y,
                                          input_state.user_inputs.diamond.x,
                                          input_state.user_inputs.diamond.b,
                                          input_state.user_inputs.diamond.a
                );
        }
        case access_read_dials: {
            apb_response.prdata = bundle( input_state.inputs_changed,
                                          13b0,
                                          input_state.user_inputs.right_dial.pressed,
                                          input_state.user_inputs.left_dial.pressed,
                                          input_state.right_dial_position,
                                          input_state.left_dial_position);
        }
        }

        /*b All done */
    }

    /*b Handle the input state */
    input_logic """
    The input state logic is relatively simple.

    The current @a user_inputs are recorded on @a
    input_state.user_inputs. When a change is detected, @a
    inputs_changed is asserted; this is only cleared on a read of the
    state register.

    The rotary dial's positions are updated when the @a
    direction_pulse asserts, using the appropriate @a dial_direction
    to indicate whether to increment or decrement.
    """: {
        if (access==access_read_state) {
            input_state.inputs_changed <= 0;
        }

        input_state.user_inputs <= user_inputs;
        if (input_state.user_inputs.left_dial.direction_pulse) {
            input_state.inputs_changed <= 1;
            if (input_state.user_inputs.left_dial.direction) {
                input_state.left_dial_position <= input_state.left_dial_position - 1;
            } else {
                input_state.left_dial_position <= input_state.left_dial_position + 1;
            }
        }
        if (input_state.user_inputs.right_dial.direction_pulse) {
            input_state.inputs_changed <= 1;
            if (input_state.user_inputs.right_dial.direction) {
                input_state.right_dial_position <= input_state.right_dial_position - 1;
            } else {
                input_state.right_dial_position <= input_state.right_dial_position + 1;
            }
        }
        if (user_inputs.diamond.a != input_state.user_inputs.diamond.a) { input_state.inputs_changed <= 1; }
        if (user_inputs.diamond.b != input_state.user_inputs.diamond.b) { input_state.inputs_changed <= 1; }
        if (user_inputs.diamond.x != input_state.user_inputs.diamond.x) { input_state.inputs_changed <= 1; }
        if (user_inputs.diamond.y != input_state.user_inputs.diamond.y) { input_state.inputs_changed <= 1; }
        if (user_inputs.joystick.u != input_state.user_inputs.joystick.u) { input_state.inputs_changed <= 1; }
        if (user_inputs.joystick.d != input_state.user_inputs.joystick.d) { input_state.inputs_changed <= 1; }
        if (user_inputs.joystick.l != input_state.user_inputs.joystick.l) { input_state.inputs_changed <= 1; }
        if (user_inputs.joystick.r != input_state.user_inputs.joystick.r) { input_state.inputs_changed <= 1; }
        if (user_inputs.joystick.c != input_state.user_inputs.joystick.c) { input_state.inputs_changed <= 1; }
        if (user_inputs.left_dial.pressed  != input_state.user_inputs.left_dial.pressed)  { input_state.inputs_changed <= 1; }
        if (user_inputs.right_dial.pressed != input_state.user_inputs.right_dial.pressed) { input_state.inputs_changed <= 1; }
        if (user_inputs.touchpanel_irq != input_state.user_inputs.touchpanel_irq) { input_state.inputs_changed <= 1; }
        if (user_inputs.temperature_alarm != input_state.user_inputs.temperature_alarm) { input_state.inputs_changed <= 1; }
    }

    /*b Done
     */
}

/*a Editor preferences and notes
mode: c ***
c-basic-offset: 4 ***
c-default-style: (quote ((c-mode . "k&r") (c++-mode . "k&r"))) ***
outline-regexp: "/\\\*a\\\|[\t ]*\/\\\*[b-z][\t ]" ***
*/
