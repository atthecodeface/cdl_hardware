/** Copyright (C) 2019,  Gavin J Stark.  All rights reserved.
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *   http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * @file  tb_apb_target_i2c.cdl
 * @brief Testbench for APB processor (ROM-based APB trasanctions)
 *
 * This is a simple testbench for the ROM-based APB transaction processor
 */
/*a Includes */
include "types/apb.h"
include "types/i2c.h"
include "input/i2c_modules.h"
include "apb/apb_targets.h"

/*a External modules */
extern module se_test_harness( clock clk,
                               output t_apb_request  apb_request,
                               input t_apb_response  apb_response,
                               input  t_i2c i2c_in,
                               output t_i2c i2c_out,
                               output t_i2c_conf i2c_conf,
                               input  bit[16] gpio_output
    )
{
    timing from rising clock clk apb_request, i2c_out, i2c_conf;
    timing to   rising clock clk apb_response, i2c_in, gpio_output;
}

/*a Module */
module tb_apb_target_i2c( clock clk,
                               input bit reset_n
)
{

    /*b Nets */
    net t_apb_request   apb_request;
    net t_apb_response  apb_response;
    net t_apb_request   i2c_apb_request;
    net t_apb_response  i2c_apb_response;
    comb t_i2c i2c_in;
    net t_i2c i2c_th;
    net t_i2c i2c_slave;
    net t_i2c i2c_master;

    net t_i2c_conf i2c_conf;
    comb t_i2c_slave_select slave_select;
    net t_i2c_action i2c_action;
    net t_i2c_slave_request slave_request;
    net t_i2c_slave_response slave_response;
    net bit[16] gpio_output;
    net bit[16] gpio_output_enable;

    /*b Instantiations */
    instantiations: {
        i2c_in  = i2c_th;
        // i2c_in &= i2c_slave;
        i2c_in.scl = i2c_in.scl & i2c_slave.scl;
        i2c_in.sda = i2c_in.sda & i2c_slave.sda;
        i2c_in.scl = i2c_in.scl & i2c_master.scl;
        i2c_in.sda = i2c_in.sda & i2c_master.sda;
        slave_select = {mask=7h70, value=7h10};
        se_test_harness th( clk <- clk,
                            apb_request => apb_request,
                            apb_response <= apb_response,
                            i2c_in  <= i2c_in,
                            i2c_out => i2c_th,
                            i2c_conf => i2c_conf,
                            gpio_output <= gpio_output
            );

        apb_target_i2c_master apb_i2c( clk <- clk,
                                       reset_n <= reset_n,
                                       apb_request  <= apb_request,
                                       apb_response => apb_response,
                                       i2c_in  <= i2c_in,
                                       i2c_out => i2c_master );

        i2c_interface i2c( clk <- clk,
                           reset_n <= reset_n,
                           i2c_in <= i2c_in,
                           i2c_action => i2c_action,
                           i2c_conf <= i2c_conf );
        
        i2c_slave slave(clk <- clk,
                        reset_n    <= reset_n,
                        i2c_action <= i2c_action,
                        i2c_out    => i2c_slave,
                        slave_select   <= slave_select, 
                        slave_request  => slave_request,
                        slave_response <= slave_response );

        i2c_slave_apb_master i2c_apb( clk <- clk,
                                      reset_n <= reset_n,
                                      slave_request <= slave_request,
                                      slave_response => slave_response,
                                      apb_request => i2c_apb_request,
                                      apb_response <= i2c_apb_response );
        apb_target_gpio gpio(clk <- clk,
                             reset_n <= reset_n,
                             apb_request <= i2c_apb_request,
                             apb_response => i2c_apb_response,
                             gpio_output => gpio_output,
                             gpio_output_enable => gpio_output_enable,
                             gpio_input <= gpio_output);
    }

    /*b All done */
}
