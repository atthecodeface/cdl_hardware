/** @copyright (C) 2019,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   vcu108_riscv.cdl
 * @brief  RISC-V design for the VCU108 board
 *

 */

/*a Includes
 */
include "subsystem/subsys_minimal.h"
include "types/video.h"
include "types/apb.h"
include "types/csr.h"
include "types/dprintf.h"
include "types/sram.h"
include "types/uart.h"
include "types/memories.h"
include "types/ethernet.h"
include "srams.h"
include "apb/apb_targets.h"
include "apb/apb_masters.h"
include "csr/csr_targets.h"
include "csr/csr_masters.h"
include "utils/dprintf_modules.h"
include "utils/async_reduce_modules.h"
include "led/led_modules.h"
include "video/framebuffer_modules.h"
include "networking/ethernet_modules.h"
include "networking/gmii_modules.h"
include "cpu/riscv/riscv_modules.h"
include "boards/vcu108.h"

typedef bit[32] t_bit32;

/*a Constants */
constant integer num_dprintf_requesters=4;

/*a Module
 */
/*m vcu108_riscv
 *
 * Debug module for testing out HPS in the Cyclone-V FPGA
 *
 */
module vcu108_riscv_3( clock clk,
                     clock clk_50,
                     input bit reset_n,

                     input  t_dprintf_req_4 vcu108_dprintf_req "Dprintf request from board (sync to clk)",
                     output bit             vcu108_dprintf_ack "Ack for dprintf request",
                     input  t_vcu108_inputs vcu108_inputs,
                     output t_vcu108_outputs vcu108_outputs,

                     clock video_clk,
                     input bit video_reset_n,
                     output t_adv7511 vcu108_video,

                     clock     sgmii_tx_clk       "Four-bit transmit serializing data clock (312.5MHz)",
                     input bit sgmii_tx_reset_n   "Reset deasserting sync to sgmii_tx_clk",
                     output bit[4] sgmii_txd      "First bit for wire in txd[0]",

                     clock     sgmii_rx_clk       "Four-bit receive serializing data clock (312.5MHz)",
                     input bit sgmii_rx_reset_n   "Reset deasserting sync to sgmii_rx_clk",
                     input bit[4] sgmii_rxd       "Oldest bit in rxd[0]",
                     output  t_sgmii_transceiver_control sgmii_transceiver_control  "Control of transceiver, on sgmii_rx_clk",
                     input t_sgmii_transceiver_status    sgmii_transceiver_status   "Status from transceiver, on sgmii_rx_clk",

                     clock flash_clk,
                     input t_mem_flash_in flash_in,
                     output t_mem_flash_out flash_out
    )
{
    /*b Clock and reset */
    default clock clk;
    default reset active_low reset_n;

    /*b Nets */
    net  t_apb_request riscv_apb_request;
    net t_apb_response riscv_apb_response;

    comb t_apb_request rv_sram_apb_request;
    comb t_apb_request riscv_dbg_apb_request;

    net t_apb_response  rv_sram_apb_response;
    net t_apb_response  riscv_dbg_apb_response;

    net t_timer_control timer_control;
    net bit[32] rv_sram_ctrl;

    net bit[num_dprintf_requesters]                 dprintf_ack;
    clocked t_dprintf_req_4[num_dprintf_requesters] dprintf_req={*=0};
    net bit[num_dprintf_requesters-1]               mux_dprintf_ack "Ack for dprintf request after multiplexing";
    net t_dprintf_req_4[num_dprintf_requesters-1]   mux_dprintf_req "Dprintf request after multiplexing";

    net bit                                         fifo_dprintf_ack "Ack for dprintf request after multiplexing";
    net t_dprintf_req_4                             fifo_dprintf_req "Dprintf request after multiplexing";

    net t_video_bus video_bus;

    net  t_riscv_debug_mst   riscv_debug_mst;
    net t_riscv_debug_tgt    riscv_debug_tgt;
    comb t_riscv_config riscv_config;
    net t_riscv_i32_trace riscv_trace;
    comb t_riscv_irqs       irqs;
    net t_sram_access_req  rv_sram_access_req;
    net t_sram_access_resp rv_sram_access_resp;

    net t_axi4s32 rx_axi4s;
    net bit       rx_axi4s_tready;
    net t_axi4s32 tx_axi4s;
    net bit       tx_axi4s_tready;
    comb t_tbi_valid tbi_rx;
    net bit[4] sgmii_txd_r;
    net bit gmii_rx_enable;
    net t_gmii_rx gmii_rx;
    net t_gmii_tx gmii_tx;
    net bit gmii_tx_enable;
    clocked t_sgmii_gasket_control sgmii_gasket_control = {*=0};
    net t_sgmii_gasket_status sgmii_gasket_status;
    clocked bit eth_reset_n = 0;

    clocked bit[32] analyzer_mux_control=0;
    clocked bit[32] analyzer_trace = {*=0};
    clocked t_bit32[8] traces = {*=0};
    
    clocked t_vcu108_inputs vcu108_inputs_r = {*=0};
    clocked bit[16] counter=0;
    clocked bit last_second_toggle=0;
    clocked bit divider_reset=0;
    clocked bit[32][4] per_sec_counters={*=0};

    default clock clk_50;
    clocked bit[32] divider=0;
    clocked bit     second_toggle=0;
    clocked bit[8]  seconds=0;

    default clock video_clk;
    default reset active_low video_reset_n;
    clocked t_adv7511 vcu108_video={*=0};
    clocked bit[4] vga_seconds_sr = 0;
    clocked bit[32][4] vga_counters={*=0};

    default clock flash_clk;
    default reset active_low reset_n;
    clocked t_mem_flash_out flash_out={*=0};

    /*b Subsystem */
    net t_csr_request   csr_request;
    net t_csr_response  csr_response;
    comb  t_subsys_inputs   subsys_inputs;
    net t_subsys_outputs  subsys_outputs;
    subsystem_instance : {
        subsys_inputs = {*=0};
        subsys_inputs.i2c = vcu108_inputs.i2c;
        subsys_inputs.uart_rx  = vcu108_inputs.uart_rx;
        subsys_inputs.switches[4;0] = vcu108_inputs.switches;
        analyzer_mux_control <= 0;
        vcu108_outputs.i2c     = subsys_outputs.i2c;
        vcu108_outputs.uart_tx = subsys_outputs.uart_tx;
        subsys_minimal subsys( clk <- clk,
                               reset_n <= reset_n,

                               master_apb_request <= riscv_apb_request,
                               master_apb_response => riscv_apb_response,

                               master_dprintf_req <= fifo_dprintf_req,
                               master_dprintf_ack => fifo_dprintf_ack,

                               master_csr_request  => csr_request,
                               master_csr_response <= csr_response,

                               subsys_inputs <= subsys_inputs,
                               subsys_outputs => subsys_outputs,

                               video_clk     <- video_clk,
                               video_reset_n <= video_reset_n,
                               
                               video_bus => video_bus,
                               tx_axi4s_tready <= tx_axi4s_tready,
                               tx_axi4s => tx_axi4s,
                               rx_axi4s <= rx_axi4s,
                               rx_axi4s_tready => rx_axi4s_tready,
                               timer_control => timer_control,
                               analyzer_trace <= analyzer_trace
            );
    }
    
    /*b RISC-V */
    riscv_instance: {
        riscv_config = {*=0};
        riscv_config.e32   = 0;
        riscv_config.i32c  = 1;
        irqs = {*=0};
        // irqs.mtip = timer_value.irq;
        riscv_i32_minimal3 riscv(clk     <- clk,
                                 proc_reset_n <= reset_n & rv_sram_ctrl[0],
                                 reset_n <= reset_n,
                                 irqs         <= irqs,
                                 sram_access_req <= rv_sram_access_req,
                                 sram_access_resp => rv_sram_access_resp,
                                      apb_request  => riscv_apb_request,
                                      apb_response <= riscv_apb_response,
                                 debug_mst <= riscv_debug_mst,
                                 debug_tgt =>riscv_debug_tgt,
                                 riscv_config <= riscv_config,
                                 trace => riscv_trace
            );
        riscv_i32_trace trace(clk <- clk,
                              reset_n <= reset_n,
                              riscv_clk_enable <= 1,
                              trace <= riscv_trace );
        riscv_i32_debug rv_debug( clk <- clk, reset_n <= reset_n,
                                  apb_request  <= riscv_dbg_apb_request,
                                  apb_response =>  riscv_dbg_apb_response,

                                  debug_mst => riscv_debug_mst,
                                  debug_tgt <= riscv_debug_tgt );
    }

    /*b Dprintf requesting */
    dprintf_requesting : {
        for (i; num_dprintf_requesters) {
            if (dprintf_ack[i]) {
                dprintf_req[i].valid <= 0;
            }
        }
        if (divider_reset) {
            dprintf_req[1] <= {valid=1, address=440,
                    data_0=bundle(32h56_47_41_3a, 32h_00_00_00_87), // VGA:%08x %08x %08x (cnts0/1/2)
                    data_1=bundle(vga_counters[0], 32h20000087),
                    data_2=bundle(vga_counters[1], 32h20000087),
                    data_3=bundle(vga_counters[2], 8hff, 24h0) };
        }
        if (divider_reset) {
            dprintf_req[0] <= {valid=1, address=400,
                    data_0=bundle(32h44_49_56_3a, 32h_00_00_00_87), // DIV:%08x %08x %08x (cnts0/1/2)
                    data_1=bundle(per_sec_counters[0], 32h20000087),
                    data_2=bundle(per_sec_counters[1], 32h20000087),
                    data_3=bundle(per_sec_counters[2], 8hff, 24h0) };
        }

        vcu108_dprintf_ack = 1;
        if (dprintf_req[2].valid) {
            vcu108_dprintf_ack = 0;
            if (dprintf_ack[2]) {
                dprintf_req[2].valid <= 0;
            }
        } else {
            if (vcu108_dprintf_req.valid) {
                dprintf_req[2] <= vcu108_dprintf_req;
            }
        }

        for (i; num_dprintf_requesters) {
            if (rv_sram_ctrl[24+i]) {
                dprintf_req[i].valid <= 0;
            }
        }
    }

    /*b Dprintf multiplexing */
    dprintf_multiplexing """
    mux[n-2] = req[n-2] * req[n-1]
    mux[n-3] = req[n-2] * mux[n-2]
    mux[2]   = req[2] * mux[3]
    mux[1]   = req[1] * mux[2]
    mux[0]   = req[0] * mux[1]
    """: {
        dprintf_4_mux tdm_n( clk <- clk,
                             reset_n <= reset_n,
                             req_a <= dprintf_req[num_dprintf_requesters-2],
                             ack_a => dprintf_ack[num_dprintf_requesters-2],
                             req_b <= dprintf_req[num_dprintf_requesters-1],
                             ack_b => dprintf_ack[num_dprintf_requesters-1],
                             req => mux_dprintf_req[num_dprintf_requesters-2],
                             ack <= mux_dprintf_ack[num_dprintf_requesters-2] );

        for (i; num_dprintf_requesters-2) {
            dprintf_4_mux tdm[i]( clk <- clk, reset_n <= reset_n,
                                  req_a <= dprintf_req[i],
                                  ack_a => dprintf_ack[i],
                                  req_b <= mux_dprintf_req[i+1],
                                  ack_b => mux_dprintf_ack[i+1],
                                  req => mux_dprintf_req[i],
                                  ack <= mux_dprintf_ack[i] );
        }
        dprintf_4_fifo_4 dpf( clk <- clk, reset_n <= reset_n,
                            req_in <= mux_dprintf_req[0],
                            ack_in => mux_dprintf_ack[0],
                            req_out => fifo_dprintf_req,
                            ack_out <= fifo_dprintf_ack );

    }

    /*b APB targets */
    comb bit[4] apb_request_sel;
    net  t_apb_request apb_request;
    comb t_apb_response apb_response;
    apb_target_instances: {
        csr_target_apb csr2apb(clk <- clk, reset_n <= reset_n,
                               csr_request  <= csr_request,
                               csr_response => csr_response,
                               apb_request  => apb_request, // top at address 0; address[16;0] from csr_request address
                               apb_response <= apb_response,
                               csr_select   <= 16h8 // csr_select field must match this
            );

        apb_request_sel = apb_request.paddr[4;10]; // in subsys_minimal 16kW
        rv_sram_apb_request           = apb_request;
        rv_sram_apb_request.psel      = apb_request.psel && (apb_request_sel==0);

        riscv_dbg_apb_request         = apb_request;
        riscv_dbg_apb_request.psel    = apb_request.psel && (apb_request_sel==1);
        
        apb_response = {*=0, pready=1};
        if (apb_request_sel==0) { apb_response = rv_sram_apb_response; }
        if (apb_request_sel==1) { apb_response = riscv_dbg_apb_response; }

        apb_target_sram_interface rv_sram_if( clk <- clk,
                                           reset_n <= reset_n,
                                           apb_request  <= rv_sram_apb_request,
                                           apb_response => rv_sram_apb_response,
                                           sram_ctrl    => rv_sram_ctrl,
                                           sram_access_req => rv_sram_access_req,
                                           sram_access_resp <= rv_sram_access_resp );

    }

    /*b Dprintf/framebuffer */
    dprintf_framebuffer_instances: {

        vcu108_video.hsync    <= video_bus.hs;
        vcu108_video.vsync    <= video_bus.vs;
        vcu108_video.de       <= video_bus.display_enable;
        vcu108_video.data[8;0]   <= video_bus.red  [8;0];
        vcu108_video.data[8;8]   <= video_bus.green[8;0];
        vcu108_video.spdif <= 0;
        //  hdmi.blue    <= bundle(video_bus.blue [8;0],2b0);

        if (video_bus.vsync) {
            vga_counters[0] <= vga_counters[0]+1;
        }
        if (video_bus.hsync) {
            vga_counters[1] <= vga_counters[1]+1;
        }
        if (video_bus.display_enable) {
            vga_counters[2] <= vga_counters[2]+1;
        }
        vga_seconds_sr <= bundle(seconds[0], vga_seconds_sr[3;1]);
        if (vga_seconds_sr[0]!=vga_seconds_sr[1]) {
            vga_counters[0] <= 0;
            vga_counters[1] <= 0;
            vga_counters[2] <= 0;
            vga_counters[3] <= 0;
        }

    }

    /*b Ethernet */
    net t_packet_stat tx_packet_stat;
    net t_packet_stat rx_packet_stat;
    ethernet : {
        gbe_axi4s32 gbe( tx_aclk <- clk,
                         tx_areset_n <= reset_n,
                         tx_axi4s    <= tx_axi4s,
                         tx_axi4s_tready => tx_axi4s_tready,
                         gmii_tx_enable <= gmii_tx_enable,
                         gmii_tx        => gmii_tx,

                         tx_packet_stat      => tx_packet_stat,
                         tx_packet_stat_ack  <= 1,

                         rx_aclk     <- clk,
                         rx_areset_n <= reset_n,
                         rx_axi4s    => rx_axi4s,
                         rx_axi4s_tready <= rx_axi4s_tready,
                         gmii_rx_enable <= gmii_rx_enable,
                         gmii_rx <= gmii_rx,

                         rx_packet_stat      => rx_packet_stat,
                         rx_packet_stat_ack  <= 1,
                         
                         rx_timer_control  <= timer_control // rx clock domain
            );

        sgmii_gasket_control.write_config  <= rv_sram_ctrl[3];
        sgmii_gasket_control.write_address <= rv_sram_ctrl[4;4];
        sgmii_gasket_control.write_data    <= bundle(8b0,rv_sram_ctrl[24;8]);
        sgmii_gmii_gasket sgg(tx_clk       <- clk,
                              tx_reset_n   <= reset_n,
                              tx_clk_312_5     <- sgmii_tx_clk,
                              tx_reset_312_5_n <= sgmii_tx_reset_n,

                              rx_clk       <- clk,
                              rx_reset_n   <= reset_n,
                              rx_clk_312_5     <- sgmii_rx_clk,
                              rx_reset_312_5_n <= sgmii_rx_reset_n,
                              
                              gmii_tx <= gmii_tx,
                              gmii_tx_enable => gmii_tx_enable,
                              // tbi_tx => tbi_tx,
                              sgmii_txd => sgmii_txd_r,

                              sgmii_rxd <= bundle(sgmii_rxd[0],sgmii_rxd[1],sgmii_rxd[2],sgmii_rxd[3]),
                              tbi_rx <= tbi_rx,
                              gmii_rx => gmii_rx,
                              gmii_rx_enable => gmii_rx_enable,
                              sgmii_gasket_control <= sgmii_gasket_control,
                              sgmii_gasket_status  => sgmii_gasket_status
            );
        tbi_rx = {*=0};
        sgmii_txd = bundle(sgmii_txd_r[0], sgmii_txd_r[1], sgmii_txd_r[2], sgmii_txd_r[3]);
    }
    
    /*b Analyzer trace */
    net bit     trace_sgmii_txd_valid;
    net bit[28] trace_sgmii_txd;
    net bit     trace_sgmii_rxd_valid;
    net bit[28] trace_sgmii_rxd;
    analyzer_trace : {
        async_reduce2_4_28_r sgmii_rxd_trace_reduce( clk_in <- sgmii_rx_clk,
                                                    clk_out <- clk,
                                                    reset_n <= reset_n,
                                                    valid_in <= 1,
                                                    data_in <= bundle(sgmii_rxd[0],sgmii_rxd[1],sgmii_rxd[2],sgmii_rxd[3]),
                                                    valid_out => trace_sgmii_rxd_valid,
                                                    data_out  => trace_sgmii_rxd );
        async_reduce2_4_28_r sgmii_txd_trace_reduce( clk_in <- sgmii_tx_clk,
                                                    clk_out <- clk,
                                                    reset_n <= reset_n,
                                                    valid_in <= 1,
                                                    data_in <= bundle(sgmii_txd[0],sgmii_txd[1],sgmii_txd[2],sgmii_txd[3]),
                                                    valid_out => trace_sgmii_txd_valid,
                                                    data_out  => trace_sgmii_txd );
        
        traces[0] <= bundle( tx_axi4s.t.data[16;0], tx_axi4s.t.user[12;0], 1b0, tx_axi4s.t.last, tx_axi4s.valid, tx_axi4s_tready );
        traces[1] <= bundle( rx_axi4s.t.data[16;0], rx_axi4s.t.user[12;0], 1b0, rx_axi4s.t.last, rx_axi4s.valid, rx_axi4s_tready );
        traces[2] <= bundle( 4b0, gmii_tx.txd, 1b0, gmii_tx.tx_er, gmii_tx.tx_en, gmii_tx_enable,
                             4b0, gmii_rx.rxd, gmii_rx.rx_crs, gmii_rx.rx_er, gmii_rx.rx_dv, gmii_rx_enable );
        traces[3] <= sgmii_gasket_status.an_state;
        traces[4] <= bundle( sgmii_gasket_status.rx_symbols_since_sync[24;0], 6b0, sgmii_gasket_status.rx_sync_toggle, sgmii_gasket_status.rx_sync);
        traces[5] <= bundle( trace_sgmii_txd, 3b0, trace_sgmii_txd_valid);
        traces[6] <= bundle( trace_sgmii_rxd, 3b0, trace_sgmii_rxd_valid);
        analyzer_trace <= traces[0];
        full_switch (analyzer_mux_control) {
        case 0: { analyzer_trace <= traces[0]; }
        case 1: { analyzer_trace <= traces[1]; }
        case 2: { analyzer_trace <= traces[2]; }
        case 3: { analyzer_trace <= traces[3]; }
        case 4: { analyzer_trace <= traces[4]; }
        case 5: { analyzer_trace <= traces[5]; }
        case 6: { analyzer_trace <= traces[6]; }
        case 7: { analyzer_trace <= traces[7]; }
        default: { analyzer_trace <= traces[0]; }
        }
    }
    /*b Second divider and second_toggle - on clk_50MHz which won't change frequency */
    second_divider : {
        /*b 50MHz stuff */
        divider <= divider+1;
        if (divider==50*1000*1000) {
            divider <= 0;
            second_toggle <= !second_toggle;
            seconds <= seconds + 1;
        }
    }

    /*b SGMII RX clock domain debug */
    default clock sgmii_rx_clk;
    default reset active_low sgmii_rx_reset_n;
    clocked bit[64] sgmii_sr = 0;
    clocked bit[64] sgmii_data = 0;
    clocked bit[8] sgmii_divider_reset_delay = 0;
    sgmii_rx_debug : {
        sgmii_sr       <= sgmii_sr>>4;
        sgmii_sr[4;60] <= sgmii_rxd;

        if (sgmii_divider_reset_delay[0]) { // Capture data for display a number of clock ticks after reset so it is stable
            full_switch (vcu108_inputs.switches[2;1]) {
            case 0: { sgmii_data <= sgmii_sr; }
            case 1: { sgmii_data <= sgmii_sr; }
            case 2: { sgmii_data <= sgmii_sr; }
            case 3: { sgmii_data <= sgmii_sr; }
            }
        }
        sgmii_divider_reset_delay <= sgmii_divider_reset_delay>>1;
        sgmii_divider_reset_delay[7] <= divider_reset;
    }
    
    /*b Stub out unused outputs and all done */
    stubs : {
        if (!sgmii_gasket_status.rx_sync) { per_sec_counters[0] <= per_sec_counters[0] + (32h1<<28); }
        per_sec_counters[0][16;0]  <= sgmii_gasket_status.an_config;
        per_sec_counters[0][12;16] <= sgmii_gasket_status.an_state[12;0];
        per_sec_counters[1] <= sgmii_data[32;0];
        per_sec_counters[2] <= sgmii_data[32;32];
            
        /*b Clock stuff */
        last_second_toggle <= second_toggle;
        divider_reset <= 0;
        if (last_second_toggle!=second_toggle) {
            divider_reset <= 1;
        }
        if (divider_reset) {
            for (i; 4) {
                per_sec_counters[i] <= 0;
            }
        }

        vcu108_inputs_r <= vcu108_inputs;        
        full_switch (vcu108_inputs.switches[2;1]) {
        case 0: { if (mux_dprintf_req[0].valid)         { counter <= counter + 1; } }
        case 1: { if (apb_request.psel)                 { counter <= counter + 1; } }
        case 3: { if (gmii_rx_enable)                   { counter <= counter + 1; } }
        }

        vcu108_outputs.i2c_reset_mux_n = subsys_outputs.gpio_output_enable[2] ? subsys_outputs.gpio_output[2] : 1;

        flash_out <= {*=0}; // wp, reset not used
        flash_out.we_n <= 1;
        flash_out.adv_n <= 1;
        flash_out.oe_n <= 1;
        flash_out.ce_n <= 1;
        flash_out.data_enable <= 0;
        
        vcu108_outputs.mdio = { mdc=1, mdio=1, mdio_enable=0 };
        eth_reset_n <= 1; // async reset to 0
        vcu108_outputs.eth_reset_n = eth_reset_n;
        
        vcu108_outputs.leds = counter[8;0];

        sgmii_transceiver_control  = {*=0};
    }
}
