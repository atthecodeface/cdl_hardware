/** Copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *   http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * @file   picoriscv_de1_cl.cdl
 * @brief  Pico-RISC-V microcomputer for the CL DE1 + daughterboard
 *
 * CDL module containing the pico-RISC-V microcomputer for the
 * Cambridge University Computer Laboratory DE1 + daughterboard
 * system.
 *
 */
/*a Includes */
include "picoriscv_types.h"
include "picoriscv.h"
include "de1_cl.h"
include "dprintf.h"
include "input_devices.h"
include "leds.h"
include "de1_cl.h"

/*a Module */
module picoriscv_de1_cl( clock clk          "50MHz clock from DE1 clock generator",
                         clock video_clk    "9MHz clock from PLL, derived from 50MHz",
                         input bit reset_n  "hard reset from a pin - a key on DE1",
                         input bit video_locked "High if video PLL has locked",
                         output t_de1_cl_lcd lcd   "LCD display out to computer lab daughterboard",
                         input bit[4] keys       "DE1 keys",
                         input bit[10] switches  "DE1 switches",
                         output bit[10] leds     "DE1 leds",
                         input t_ps2_pins ps2_in   "PS2 input pins",
                         output t_ps2_pins ps2_out "PS2 output pin driver open collector",
                         output bit led_data_pin "DE1 CL daughterboard neopixel LED pin",
                         input  t_de1_cl_inputs_status   inputs_status  "DE1 CL daughterboard shifter register etc status",
                         output t_de1_cl_inputs_control  inputs_control "DE1 CL daughterboard shifter register control"
    )
{
    net t_video_bus prv_video_bus;
    comb t_video_bus io_video_bus;

    //net t_ps2_pins ps2_out;

    comb t_csr_request csr_request;
    net t_csr_response prv_csr_response;

    comb  bit led_chain;
    //net bit[10] leds;
    //net  t_de1_cl_inputs_control inputs_control "DE1 CL IO inputs control - shift register clock, and so on";

    comb bit prv_reset_n;
    comb bit video_reset_n;
    comb t_prv_keyboard prv_keyboard;
    comb bit lcd_source;

    /*b Miscellaneous logic */
    misc_logic """
    """: {
        prv_reset_n       = reset_n & switches[0]; // & !prv_clock_control.reset_cpu;
        video_reset_n     = reset_n & video_locked;
    }

    /*b DE1/CL IO for PRV subsystem */
    prv_de1_cl_instantiations: {
        lcd_source = 0;
        prv_keyboard = {*=0};
        led_chain = 0;
        csr_request = {*=0};
        io_video_bus = {*=0};
        inputs_control = {*=0};
        ps2_out = {*=0};
        leds = 0;
        /*
        picoriscv_de1_cl_io io( clk <- clk,
                                video_clk <- video_clk,
                                reset_n <= reset_n,
                                prv_reset_n <= prv_reset_n,
                                framebuffer_reset_n <= framebuffer_reset_n,
                                keys <= keys,
                                switches <= switches,
                                clock_control <= prv_clock_control,
                                prv_keyboard => prv_keyboard,
                                video_bus => io_video_bus,
                                csr_request => csr_request,
                                csr_response <= prv_csr_response,
                                inputs_control => inputs_control,
                                inputs_status <= inputs_status,
                                ps2_in <= ps2_in,
                                ps2_out => ps2_out,
                                lcd_source => lcd_source,
                                leds => leds,
                                led_chain => led_chain
            );
        */
    }

    /*b PRV Micro subsystem */
    picoriscv_instantiations: {
        picoriscv prv( clk <- clk,
                       video_clk <- video_clk,
                       reset_n <= prv_reset_n,
                       video_reset_n <= video_reset_n,
                       keyboard <= prv_keyboard,
                       video_bus => prv_video_bus,
                       csr_request <= csr_request,
                       csr_response => prv_csr_response );
    }

    /*b Output muxes */
    output_muxes """
    """: {
        lcd = { vsync_n        = !prv_video_bus.vsync,
                hsync_n        = !prv_video_bus.hsync,
                display_enable = prv_video_bus.display_enable,
                red            = prv_video_bus.red[6;2],
                green          = prv_video_bus.green[7;1],
                blue           = prv_video_bus.blue[6;2],
                backlight = switches[1]
        };
        if (lcd_source) {
            lcd = { vsync_n        = !io_video_bus.vsync,
                    hsync_n        = !io_video_bus.hsync,
                    display_enable = io_video_bus.display_enable,
                    red            = io_video_bus.red[6;2],
                    green          = io_video_bus.green[7;1],
                    blue           = io_video_bus.blue[6;2]
            };
        }
        led_data_pin = !led_chain;
    }

    /*b All done */
}
