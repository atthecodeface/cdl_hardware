/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   riscv_simple.cdl
 * @brief  Very simple RISC-V implementation ported to CDL
 *
 * CDL implementation of very simple RISC-V teaching implementation
 *
 */

/*a Includes
 */
include "riscv_internal_types.h"
include "riscv.h"
include "riscv_submodules.h"

/*a Constants
 */
constant integer INITIAL_PC=0x0;
constant integer i32c_force_disable=0;

/*a Types
 */
/*t t_decexec_state */
typedef struct {
    t_riscv_i32_inst instruction   "Fetched instruction, ready for decode, register fetch, execute and writeback";
    bit valid;
    bit[32] pc                   "PC of the decoded instruction";
} t_decexec_state;

/*t t_decexec_combs
 *
 * Combinatorials of the decexec_state
 */
typedef struct {
    t_riscv_i32_decode idecode;

    t_riscv_word   rs1;
    t_riscv_word   rs2;
    bit[32] next_pc;

    bit[2]  word_offset;
    bit branch_taken;
    t_riscv_csr_access csr_access;
} t_decexec_combs;

/*t t_rfw_state */
typedef struct {
    t_riscv_i32_decode idecode;
    bit valid;
    bit memory_read;
    bit[2]  word_offset;
    t_riscv_word result;
} t_rfw_state;

/*t t_rfw_combs
 * Combinatorial decode of rfw_state
 */
typedef struct {
    t_riscv_word write_data;
    t_riscv_word memory_data;
} t_rfw_combs;

/*a Module
 */
module riscv_i32c_pipeline2( clock clk,
                             input bit reset_n,
                             input t_riscv_irqs       irqs               "Interrupts in to the CPU",
                             output t_riscv_mem_access_req  dmem_access_req,
                             input  t_riscv_mem_access_resp dmem_access_resp,
                             output t_riscv_fetch_req       ifetch_req,
                             input  t_riscv_fetch_resp      ifetch_resp,
                             input  t_riscv_config          riscv_config,
                             output t_riscv_i32_trace       trace
)
"""
"""
{

    /*b State and comb
     */
    default clock clk;
    default reset active_low reset_n;

    clocked t_riscv_word[32] registers={*=0} "Register 0 is tied to 0 - so it is written on every cycle to zero...";

    net     t_riscv_i32_decode decexec_idecode_i32;
    net     t_riscv_i32_decode decexec_idecode_i32c;
    clocked t_decexec_state    decexec_state={*=0, pc=INITIAL_PC};
    comb    t_decexec_combs    decexec_combs;
    net     t_riscv_i32_alu_result decexec_alu_result;

    clocked t_rfw_state    rfw_state={*=0};
    comb    t_rfw_combs    rfw_combs;

    comb t_riscv_csr_controls csr_controls;
    net t_riscv_csr_data csr_data;

    /*b Ifetch stage
     */
    instruction_fetch_stage """
    The instruction fetch request derives from the
    decode/execute stage (the instruction address that is required
    next) and presents that to the outside world.

    This request may be for any 16-bit aligned address, and two
    successive 16-bit words from that request must be presented,
    aligned to bit 0.

    If the decode/execute stage is invalid (i.e. it does not have a
    valid instruction to decode) then the current PC is requested.
    """: {
        ifetch_req               = {*=0};
        // sequential?
        ifetch_req.valid         = 1;
        ifetch_req.address       = decexec_combs.next_pc;
        if (!decexec_state.valid) {
            ifetch_req.address   = decexec_state.pc;
        }
    }

    /*b Decode, RFR and execute stage
     */
    decode_rfr_execute_stage: {
        /*b Instruction register */
        decexec_state.valid <= 0;
        if (ifetch_req.valid && ifetch_resp.valid) {
            decexec_state.valid <= 1;
            decexec_state.instruction <= {data=ifetch_resp.data, mode=rv_mode_machine};
        }
        if (decexec_state.valid) {
            decexec_state.pc <= decexec_combs.next_pc;
        }

        /*b Decode instruction */
        riscv_i32_decode decode_i32( instruction <= decexec_state.instruction,
                                     idecode      => decexec_idecode_i32,
                                     riscv_config <= riscv_config );

        riscv_i32c_decode decode_i32c( instruction <= decexec_state.instruction,
                                       idecode      => decexec_idecode_i32c,
                                       riscv_config <= riscv_config );

        /*b Select decode */
        decexec_combs.idecode = decexec_idecode_i32;
        if ((!i32c_force_disable) && riscv_config.i32c) {
            if (decexec_state.instruction.data[2;0]!=2b11) {
                decexec_combs.idecode = decexec_idecode_i32c;
            }
        }

        /*b Register read */
        decexec_combs.rs1 = registers[decexec_combs.idecode.rs1]; // note that register 0 is ALWAYS 0 anyway
        decexec_combs.rs2 = registers[decexec_combs.idecode.rs2]; // note that register 0 is ALWAYS 0 anyway
        if (rfw_state.valid && rfw_state.idecode.rd_written) {
            if (decexec_combs.idecode.rs1 == rfw_state.idecode.rd) {decexec_combs.rs1 = rfw_combs.write_data;}
            if (decexec_combs.idecode.rs2 == rfw_state.idecode.rd) {decexec_combs.rs2 = rfw_combs.write_data;}
        }

        /*b Execute ALU stage */
        riscv_i32_alu alu( idecode <= decexec_combs.idecode,
                           pc  <= decexec_state.pc,
                           rs1 <= decexec_combs.rs1,
                           rs2 <= decexec_combs.rs2,
                           alu_result => decexec_alu_result );

        /*b Minimal CSRs */
        csr_controls = {*=0};
        csr_controls.retire      = decexec_state.valid;
        csr_controls.timer_inc   = 1;

        decexec_combs.csr_access = decexec_combs.idecode.csr_access;
        if (!decexec_state.valid || decexec_combs.idecode.illegal) {
            decexec_combs.csr_access.access = riscv_csr_access_none;
        }
        riscv_csrs_minimal csrs( clk <- clk,
                                 reset_n <= reset_n,
                                 irqs <= irqs,
                                 csr_access <= decexec_combs.csr_access,
                                 csr_data  => csr_data,
                                 csr_controls <= csr_controls );

        /*b Memory access */
        dmem_access_req.read_enable  = (decexec_combs.idecode.op == riscv_op_load);
        dmem_access_req.write_enable = (decexec_combs.idecode.op == riscv_op_store);
        dmem_access_req.address      = decexec_alu_result.arith_result;
        decexec_combs.word_offset    = decexec_alu_result.arith_result[2;0];
        dmem_access_req.byte_enable  = 4hf << decexec_combs.word_offset;
        part_switch (decexec_combs.idecode.memory_width) {
        case mw_byte: { dmem_access_req.byte_enable  = 4h1 << decexec_combs.word_offset; }
        case mw_half: { dmem_access_req.byte_enable  = 4h3 << decexec_combs.word_offset; }
        }
        dmem_access_req.write_data = decexec_combs.rs2 << (bundle(decexec_combs.word_offset,3b0));

        /*b Determine whether branch would be taken and find next PC */
        decexec_combs.branch_taken = 0;
        full_switch (decexec_combs.idecode.op) {
        case riscv_op_branch:   { decexec_combs.branch_taken = decexec_alu_result.branch_condition_met; }
        case riscv_op_jal:      { decexec_combs.branch_taken=1; }
        case riscv_op_jalr:     { decexec_combs.branch_taken=1; }
        }
        decexec_combs.next_pc = decexec_state.pc + 4;
        if (decexec_combs.branch_taken) {
            decexec_combs.next_pc = decexec_alu_result.branch_target;
        }

        /*b All done */
    }

    /*b RFW, memory complete stage
     */
    rfw_stage: {
        /*b Instruction register */
        rfw_state.valid <= 0;
        if (decexec_state.valid) {
            rfw_state.valid <= 1;
            rfw_state.idecode <= decexec_combs.idecode;
            if (decexec_combs.idecode.rd==0) {
                rfw_state.idecode.rd_written <= 0;
            }
            rfw_state.memory_read <= (decexec_combs.idecode.op==riscv_op_load);
            rfw_state.word_offset <= decexec_combs.word_offset;
            rfw_state.result      <= decexec_alu_result.result;
            if (decexec_combs.idecode.csr_access.access != riscv_csr_access_none) {
                rfw_state.result <= csr_data.read_data;
            }
        }

        rfw_combs.memory_data = dmem_access_resp.read_data;
        part_switch (rfw_state.idecode.memory_width) {
        case mw_byte: {
            rfw_combs.memory_data = (dmem_access_resp.read_data >> (bundle(rfw_state.word_offset,3b0))) & 0xff;
            if (!rfw_state.idecode.memory_read_unsigned && rfw_combs.memory_data[7]) { rfw_combs.memory_data[24;8] = -1; }
        }
        case mw_half: {
            rfw_combs.memory_data = (dmem_access_resp.read_data >> (bundle(rfw_state.word_offset,3b0))) & 0xffff;
            if (!rfw_state.idecode.memory_read_unsigned && rfw_combs.memory_data[15]) { rfw_combs.memory_data[16;16] = -1; }
        }
        }

        rfw_combs.write_data = rfw_state.memory_read ? rfw_combs.memory_data : rfw_state.result;
        if (rfw_state.valid && rfw_state.idecode.rd_written) {
            registers[rfw_state.idecode.rd] <= rfw_combs.write_data;
        }
        registers[0] <= 0; // register 0 is always zero...
    }

    /*b Logging */
    logging """
    """: {
        trace = {*=0};
        trace.instr_valid    = decexec_state.valid;
        trace.instr_pc       = decexec_state.pc;
        trace.instruction    = decexec_state.instruction;
        trace.rfw_retire     = rfw_state.valid;
        trace.rfw_data_valid = rfw_state.idecode.rd_written;
        trace.rfw_rd         = rfw_state.idecode.rd;
        trace.rfw_data       = rfw_combs.write_data;
        trace.branch_taken   = decexec_combs.branch_taken;
        trace.trap           = 0;
        trace.branch_target  = decexec_alu_result.branch_target;
    }

    /*b All done */
}

