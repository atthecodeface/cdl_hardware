/** Copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *   http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * @file  saa5050.cdl
 * @brief CDL implementation of Mullard SAA5050
 *
 * This is an implementaion of the 5050 teletext decoder chip, which
 * really was used in the BBC microcomputer as a teletext ROM with
 * teletext character interpretation to supply 3bpp color video from a
 * bytestream of video memory data.
 *
 * Currently this implementation does not support double-height
 * characters, blanking during control characters, or smoothing. The
 * teletext character ROM is implemented as an SRAM that is filled
 * through a host SRAM request bus - it is not readable.
 */
/*a Includes */
include "bbc_submodules.h"

/*a Types */
typedef bit[3] t_color;
/*t t_character_state */
typedef struct {
    bit[3] background_color;
    bit[3] foreground_color;
    bit    held_character;
    bit    flashing;
    bit    text_mode;
    bit    contiguous_graphics;
    bit    dbl_height;
    bit    hold_graphics;
} t_character_state;

/*t t_load_state */
typedef struct {
    bit last_lose;
    bit[7] character_data;
    bit character_data_toggle;
    bit[4] scanline;
    bit    end_of_scanline;
    bit    end_of_row;
    bit    end_of_field;
    bit[6] flashing_counter; // 50 fields per second, 3/4 second, max of ~40, flash on at 10
    bit    flash_on;
} t_load_state;
constant integer flashing_on_count=10;
constant integer max_flashing_count=40;

/*t t_pixel_decode */
typedef struct {
    bit new_character;
    bit end_of_scanline;
    bit end_of_row;
    bit end_of_field;
    t_character_state next_character_state;
    t_character_state current_character_state;
    bit can_be_replaced_with_hold;
    bit reset_held_graphics;
    bit[10] rom_scanline_data;
    bit[7] character_data;
    bit[12] smoothed_scanline_data;
} t_pixel_decode;

/*t t_pixel_state */
typedef struct {
    bit character_data_toggle;
    bit end_of_scanline;
    bit end_of_row;
    bit end_of_field;
    t_character_state character_state;
    bit[7] character_data;
    bit[2] hexpixel_of_character;
    bit row_contains_dbl_height;
    bit last_row_contained_dbl_height;
} t_pixel_state;

/*t t_hexpixel_state */
typedef struct {
    bit[6] pixels;
    t_character_state character_state;
} t_hexpixel_state;

/*a Module saa5050 */
module saa5050( clock clk_2MHz     "Supposedly 6MHz pixel clock (TR6), except we use 2MHz and deliver 3 pixels per tick; rising edge should be coincident with clk_1MHz edges",
                clock clk_1MHz     "Character clock, used to clock in the parallel data; real chip uses F1 and syncs to TR6; this clock RISES when F1 FALLS",
                input bit reset_n,
                input bit superimpose_n "Not implemented",
                input bit data_n "Serial data in, not implemented",
                input bit[7] data_in "Parallel data in",
                input bit dlim "clocks serial data in somehow (datasheet is dreadful...)",
                input bit glr "General line reset - can be tied to hsync - assert once per line before data comes in",
                input bit dew "Data entry window - used to determine flashing rate and resets the ROM decoders - can be tied to vsync",
                input bit crs "Character rounding select - drive high on even interlace fields to enable use of rounded character data (kinda indicates 'half line')",
                input bit bcs_n "Assert (low) to enable double-height characters (?) ",
                output bit tlc_n "Asserted (low) when double-height characters occur (?) ",
                input bit lose "Load output shift register enable - must be low before start of character data in a scanline, rising with (or one tick earlier?) the data; changes off falling F1, rising clk_1MHz",
                input bit de "Display enable",
                input bit po "Picture on",
                output bit[6] red,
                output bit[6] green,
                output bit[6] blue,
                output bit blan,
                input t_bbc_micro_sram_request host_sram_request "Write only, writes on clk_2MHz rising, acknowledge must be handled by supermodule"
       )
    /*b Documentation */
"""
Teletext characters are displayed from a 12x20 grid.
The ROM characters have two background rows, and then are displayed with 2 background pixels on the left, and then 10 pixels from the ROM
The ROM is actually 5x9, and it is doubled to 10x18
Doubling without smoothing can be achieved be true doubling
Doubling with smoothing is done on intervening lines:

The ROM A is:
..*..
.*.*.
*...*
*...*
*****
*...*
*...*
.....
.....

So a non-smoothed A is
....**....
....**....
..**..**..
..**..**..
**......**
**......**
**......**
**......**
**********
**********
**......**
**......**
**......**
**......**
..........
..........
..........
..........

..*..
.*.*.
*...*
*...*
*****
*...*
*...*
.....
.....

The smoothing is only to smoothe diagonals.
So the centroids are added on diagonals (baseline requirement...)
In fact, one can add 2x2 blobs on the diagonals:

A smoothed A is then:
....**....
...****...
..******..
.***..***.
***....***
**......**
**......**
**......**
**********
**********
**......**
**......**
**......**
**......**
..........
..........
..........
..........


Graphics characters are 6 blobs on a 6x10 grid (contiguous, separated):
000111 .00.11
000111 .00.11
000111 ......
222333 .22.33
222333 .22.33
222333 .22.33
222333 ......
444555 .44.55
444555 .44.55
444555 ......

The BBC micro seems to use 19 rows per character, but in practice (since it is interlaced sync and video) it will use 10 in each field, and CRS will be set for even fields


"""
{
    /*b Defaults */
    default reset active_low reset_n;
    default clock clk_1MHz;
    clocked t_load_state load_state = {*=0};
    net bit[64] pixel_rom_data;

    default clock clk_2MHz;
    clocked t_pixel_state pixel_state = {*=0};
    comb    t_pixel_decode pixel;
    clocked t_hexpixel_state hexpixel_state={*=0};
    comb t_color[6] hexpixel_colors;

    /*b Timing control and load_state stage (1MHz clock in) - scanline and character loading  */
    scanline_and_loading """
    """: {
        load_state.last_lose <= lose;
        if (lose) {
            load_state.character_data <= data_in;
            load_state.character_data_toggle <= !load_state.character_data_toggle; // change on this indicates new character to other clock
        }
        load_state.end_of_scanline <= 0;
        if (load_state.last_lose && !lose) {
            load_state.character_data <= 0;
            load_state.character_data_toggle <= !load_state.character_data_toggle; // change on this indicates new character to other clock
            load_state.scanline <= load_state.scanline+1;
            load_state.end_of_scanline <= 1;
            if (load_state.scanline==9) {
                load_state.end_of_row <= 1;
            }
        }
        if (dew) {
            load_state.end_of_row <= 1;
            load_state.end_of_field <= 1;
        }
        if (load_state.end_of_row) {
            load_state.scanline <= 0;
            load_state.character_data_toggle <= 0;
            load_state.end_of_row <= 0;
        }
        if (load_state.end_of_field) {
            load_state.flashing_counter <= load_state.flashing_counter+1;
            if (load_state.flashing_counter==flashing_on_count) {
                load_state.flash_on <= 1;
            }
            if (load_state.flashing_counter==max_flashing_count) {
                load_state.flashing_counter <= 0;
                load_state.flash_on <= 0;
            }
            load_state.end_of_field <= 0;
        }
    }

    /*b Character ROM fetch and control decode - after ROM, all is in pixel_state pipeline stage */
    character_rom_and_control_decode """
    """: {
        /*b Decode 'character_data' and scanline_of_character in ROM to get 2 lines of character
        address for ROM is character_data, and we read out 45 bits (5*9).
        Select appropriate ten bits using scanline_of_character */
        se_sram_srw_128x64 character_rom(sram_clock <- clk_2MHz,
                                         select <= 1,
                                         read_not_write <= !host_sram_request.write_enable,
                                         write_enable   <= host_sram_request.write_enable&&(host_sram_request.select==bbc_sram_select_cpu_teletext),
                                         address        <= (host_sram_request.valid&&(host_sram_request.select==bbc_sram_select_cpu_teletext)) ? host_sram_request.address[7;0] : load_state.character_data,
                                         write_data     <= host_sram_request.write_data,
                                         data_out       => pixel_rom_data );

        /*b Decode current character
          note that steady, normal size, conceal, contiguous, separated, black background, new background, hold are 'set-at'
          rest are 'set-after'.
          'set-at' means it takes immediate effect for this character, 'set-after' just for the following characters
         */
        pixel.next_character_state    = pixel_state.character_state;
        pixel.current_character_state = pixel_state.character_state;
        pixel.can_be_replaced_with_hold = 1;
        pixel.reset_held_graphics = 0;
        part_switch (load_state.character_data) {
        case 0: { // probably also the other un-interpreted <32 characters...
            pixel.can_be_replaced_with_hold = 1;
        }
        case 1,2,3,4,5,6,7: {
            pixel.next_character_state.foreground_color = load_state.character_data[3;0];
            pixel.next_character_state.text_mode = 1;
        }
        case 8: { pixel.next_character_state.flashing = 1; }
        case 9: { // steady is set-at
            pixel.current_character_state.flashing = 0;
            pixel.next_character_state.flashing = 0;
            // does this reset the held graphics?
        }
        case 17,18,19,20,21,22,23: {
            pixel.next_character_state.foreground_color = load_state.character_data[3;0];
            pixel.next_character_state.text_mode = 0;
            // does this reset the held graphics?
        }
        case 12: { // normal size is set-at
            pixel.current_character_state.dbl_height = 0;
            pixel.next_character_state.dbl_height    = 0;
            // does this reset the held graphics?
        }
        case 13: { // double height is set-after
            pixel.next_character_state.dbl_height = 1;
            // does this reset the held graphics?
        } 
        case 25: { // contiguous graphics is set-at
            pixel.current_character_state.contiguous_graphics = 1;
            pixel.next_character_state.contiguous_graphics = 1;
        }
        case 26: { // separated graphics is set-at
            pixel.current_character_state.contiguous_graphics = 0;
            pixel.next_character_state.contiguous_graphics = 0;
        }
        case 28: { // black background is set-at
            pixel.current_character_state.background_color = 0;
            pixel.next_character_state.background_color = 0;
        }
        case 29: { // new background is set-at
            pixel.current_character_state.background_color = pixel_state.character_state.foreground_color;
            pixel.next_character_state.background_color    = pixel_state.character_state.foreground_color;
        }
        case 30: { // hold mode is set-at
            pixel.next_character_state.hold_graphics = 1; // note that a held character is the last graphics character INCLUDING separated or not
            pixel.next_character_state.hold_graphics = 1;
        }
        case 31: { // release graphics is set-after
            pixel.next_character_state.hold_graphics = 0;
        }
        default: {
            pixel.can_be_replaced_with_hold = 0;
        }
        }

        /*b Handle change of control state at end of character */
        pixel_state.character_data        <= load_state.character_data;
        pixel_state.character_data_toggle <= load_state.character_data_toggle;
        pixel_state.end_of_scanline       <= load_state.end_of_scanline;
        pixel_state.end_of_row            <= load_state.end_of_row;
        pixel_state.end_of_field          <= load_state.end_of_field;
        pixel.new_character   = (pixel_state.character_data_toggle != load_state.character_data_toggle);
        pixel.end_of_scanline = (!pixel_state.end_of_scanline && load_state.end_of_scanline);
        pixel.end_of_row      = (!pixel_state.end_of_row      && load_state.end_of_row);
        pixel.end_of_field    = (!pixel_state.end_of_field    && load_state.end_of_field);

        pixel_state.hexpixel_of_character <= pixel_state.hexpixel_of_character + 1;
        if (pixel.new_character) {
            pixel_state.character_state <= pixel.next_character_state;
            pixel_state.hexpixel_of_character <= 0;
            if (pixel.current_character_state.dbl_height) {
                pixel_state.row_contains_dbl_height <= 1;
            }
        }

        /*b Handle reset of control state at end of scanline */
        if (pixel.end_of_scanline) {
            pixel_state.character_state.background_color <= 0;
            pixel_state.character_state.foreground_color <= 3b111;
            pixel_state.character_state.held_character <= 0;
            pixel_state.character_state.flashing <= 0;
            pixel_state.character_state.text_mode <= 1;
            pixel_state.character_state.contiguous_graphics <= 1;
        }

        /*b Handle reset of control state at end of character row */
        if (pixel.end_of_row) {
            pixel_state.last_row_contained_dbl_height <= pixel_state.row_contains_dbl_height;
            pixel_state.row_contains_dbl_height <= 0;
        }

        /*b Handle reset of control state at end of field */
        if (pixel.end_of_field) {
            pixel_state.last_row_contained_dbl_height <= 0;
            pixel_state.row_contains_dbl_height <= 0;
        }
    }

    /*b Character pixel generation, in pixel pipeline stage, depending on pixel.current_character_state, generating hexpixel state */
    character_pixel_generation """
    Get two scanlines - current and next (next of 0 if none)
    """: {

        /*b Select scanline of ROM data for pixel */
        full_switch (load_state.scanline) { //scanline_of_character changes every scanline, so no need to have a pixel pipeline stage version
        case 0: { pixel.rom_scanline_data = bundle(pixel_rom_data[5;0],5b0); }
        case 1: { pixel.rom_scanline_data = pixel_rom_data[10;0]; }
        case 2: { pixel.rom_scanline_data = pixel_rom_data[10;5]; }
        case 3: { pixel.rom_scanline_data = pixel_rom_data[10;10]; }
        case 4: { pixel.rom_scanline_data = pixel_rom_data[10;15]; }
        case 5: { pixel.rom_scanline_data = pixel_rom_data[10;20]; }
        case 6: { pixel.rom_scanline_data = pixel_rom_data[10;25]; }
        case 7: { pixel.rom_scanline_data = pixel_rom_data[10;30]; }
        case 8: { pixel.rom_scanline_data = pixel_rom_data[10;35]; }
        default: { pixel.rom_scanline_data = bundle(5b0,pixel_rom_data[5;35]); }
        }

        /*b Smoothe ROM data for pixel */
        // For smoothing, should smoothe if crs is set only, and text only too
        pixel.smoothed_scanline_data = bundle( 2b0,
                                               pixel.rom_scanline_data[4],pixel.rom_scanline_data[4],
                                               pixel.rom_scanline_data[3],pixel.rom_scanline_data[3],
                                               pixel.rom_scanline_data[2],pixel.rom_scanline_data[2],
                                               pixel.rom_scanline_data[1],pixel.rom_scanline_data[1],
                                               pixel.rom_scanline_data[0],pixel.rom_scanline_data[0] );

        /*b Override if in graphics mode */
        pixel.character_data = pixel_state.character_data;
        if (!pixel.current_character_state.text_mode) {
            if ((load_state.scanline==0) || (load_state.scanline==1) || (load_state.scanline==2)) {
                pixel.smoothed_scanline_data = (pixel.character_data[0]?12hfc0:12h0) | (pixel.character_data[1]?12h03f:12h0);
            } elsif ((load_state.scanline==7) || (load_state.scanline==8) || (load_state.scanline==9)) {
                pixel.smoothed_scanline_data = (pixel.character_data[4]?12hfc0:12h0) | (pixel.character_data[6]?12h03f:12h0);
            } else {
                pixel.smoothed_scanline_data = (pixel.character_data[2]?12hfc0:12h0) | (pixel.character_data[3]?12h03f:12h0);
            }
            if (!pixel.current_character_state.contiguous_graphics) {
                pixel.smoothed_scanline_data[2;10] = 2b00;
                pixel.smoothed_scanline_data[2;4]  = 2b00;
                if ((load_state.scanline==2) || (load_state.scanline==6) || (load_state.scanline==9)) {
                    pixel.smoothed_scanline_data = 0;
                }
            }
        }

        /*b Generate hexpixel_state.pixels */
        hexpixel_state.pixels <= pixel.smoothed_scanline_data[6;0];
        part_switch (pixel_state.hexpixel_of_character) {
        case 0: {hexpixel_state.pixels <= pixel.smoothed_scanline_data[6;6];}
        case 1: {hexpixel_state.pixels <= pixel.smoothed_scanline_data[6;0];}
        }
        hexpixel_state.character_state <= pixel.current_character_state;
    }

    /*b Outputs from hexpixel pipeline stage */
    outputs_from_hexpixel """
    """: {
        red = 0;
        blue = 0;
        green = 0;
        for (i; 6) {
            hexpixel_colors[i] = hexpixel_state.pixels[i] ? hexpixel_state.character_state.foreground_color : hexpixel_state.character_state.background_color;
        }
        for (i; 6) {
            red[i]   = hexpixel_colors[i][0];
            green[i] = hexpixel_colors[i][1];
            blue[i]  = hexpixel_colors[i][2];
        }
        blan = 0;
        tlc_n = 0;
    }

    /*b All done */
}
