/** @copyright (C) 2020,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   analyzer_mux_8_2e
 * @brief  Two-enabled port of analyzer_mux_8
 *
 * Needs to be built in CDL with the options:
 *
 *  dc:analyzer_config_num_targets=2
 *  rmn:analyzer_mux_8=analyzer_mux_8_e2
 *
 */
/*a Module */
include "analyzer_mux_8.cdl"
