/** Copyright (C) 2019,  Gavin J Stark.  All rights reserved.
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *   http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * @file  tb_de1_hps_generic.cdl
 * @brief Generic testbench for DE1 HPS
 *
 */
/*a Includes */
include "boards/vcu108.h"
include "boards/vcu108/vcu108_generic.h"

/*a Modules */
/*m extern for se_test_harness with extra connections */
extern
module se_test_harness(clock clk,
                       input bit reset_n,
                       output t_vcu108_inputs vcu108_inputs,
                       input t_vcu108_leds  vcu108_leds,
                       input t_adv7511 vcu108_video,
                       output bit uart_rxd,
                       input bit uart_txd
    )
{
    timing from rising clock clk vcu108_inputs, uart_rxd;
    timing to   rising clock clk vcu108_leds, vcu108_video, uart_txd;
}

/*m tb_vcu108_generic */
module tb_vcu108_generic( clock clk,
                          clock video_clk,
                          input bit reset_n
)
{

    /*b Nets */
    net t_vcu108_inputs vcu108_inputs;
    net t_vcu108_leds  vcu108_leds;

    net t_adv7511 vcu108_video;

    net bit uart_rxd;
    net bit uart_txd;

    /*b Instantiations */
    instantiations: {
        se_test_harness th(  clk <- clk,
                             reset_n <= reset_n,

                             vcu108_inputs => vcu108_inputs,
                             vcu108_leds   <= vcu108_leds,

                             vcu108_video <= vcu108_video,

                             uart_rxd => uart_rxd,
                             uart_txd <= uart_txd
            );
        
        vcu108_generic dut(  clk <- clk,
                             reset_n <= reset_n,

                             vcu108_inputs <= vcu108_inputs,
                             vcu108_leds => vcu108_leds,

                             video_clk <- video_clk,
                             video_reset_n <= reset_n,

                             vcu108_video => vcu108_video,

                             uart_rxd <= uart_rxd,
                             uart_txd => uart_txd
            );
    }

    /*b All done */
}

/*a Editor preferences and notes
mode: c ***
c-basic-offset: 4 ***
c-default-style: (quote ((c-mode . "k&r") (c++-mode . "k&r"))) ***
outline-regexp: "/\\\*a\\\|[\t ]*\/\\\*[b-z][\t ]" ***
*/
