/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   riscv_i32_decode.cdl
 * @brief  Instruction decoder for RISC-V implementation
 *
 * CDL implementation of RISC-V instruction decode based on the RISC-V
 * specification v2.2.
 *
 */

/*a Includes
 */
include "cpu/riscv/riscv_internal_types.h"
include "cpu/riscv/riscv.h"
include "cpu/riscv/riscv_config.h"
include "cpu/riscv/riscv_submodules.h"

/*a Types
 */
typedef struct {
    bit            use_debug    "Asserted if decode of instruction should be be 'debug' not regular";
    bit[2]         must_be_ones "Bits that must be one for a valid RISCV I32 base instruction";
    bit            is_imm_op "Asserted if the instruction is an immediate operation";
    bit[5]         opc     "Opcode field from 32-bit instruction";
    bit[7]         funct7  "7-bit function field of instruction";
    bit[3]         funct3  "3-bit function field of instruction";
    t_riscv_word   imm_signed "Sign-extension word, basically instruction[31] replicated";
    bit            rs1_nonzero;
} t_combs;

/*a Module
 */
module riscv_i32_decode( input t_riscv_i32_inst instruction,
                         output t_riscv_i32_decode idecode,
                         input t_riscv_config riscv_config
)
"""
Instruction decoder for RISC-V I32 instruction set.

This is based on the RISC-V v2.2 specification (hence figure numbers
are from that specification)

It provides for the option of RV32E and RV32M.

RV32E indicates an illegal instruction if a register outside 0-15 is accessed.

RV32M provides decode of multiply and divide; if it is not desired
then the instructions are decoded as illegal.

25-bit opcode spaces should chose one of the standard R/I/S/U encodings
R is Rd, Rs1, Rs2           plus 10 bits for encoding
I is Rd, Rs1, imm(12 bits)  plus 3 bits for encoding
S is Rs1, Rs2, imm(12 bits) plus 3 bits for encoding
U is Rd, imm(20 bits starting at bit 12) with no spare bits

Custom-0 is a 25-bit opcode space with instruction bottom bits of 7b0001011
Custom-1 is a 25-bit opcode space with instruction bottom bits of 7b0101011
Custom-2 is a 25-bit opcode space with instruction bottom bits of 7b1011011; this conflicts with RV-128 but is available for RV-32
Custom-3 is a 25-bit opcode space with instruction bottom bits of 7b1111011; this conflicts with RV-128 but is available for RV-32

22-bit opcode spaces are parts of the standard 25-bit opcode spaces
There are 2 unused branch encodings (funct3 of 3b010, 3b011)
There are 2 unused ALU-immediate encodings (funct3 of 3b001, 3b101)

Atomic instructions are 7b0101111 in bottom 7 bits - top 6 bits are the atomic type; this has a standard 3-register encoding

"""
{

    /*b Signals - just the combs */
    comb t_combs combs      "Combinatorials used in the module, not exported as the decode";
    comb t_riscv_i32_decode idecode_inst;
    comb t_riscv_i32_decode idecode_debug;
    comb t_riscv_csr_access csr_access "CSR access before select decode";
    net t_riscv_csr_decode  csr_decode "CSR decode (select and illegal_access) IF it were a system instruction";

    /*b Basic instruction breakout
     */
    instruction_breakout """
    Break out the instruction into fields, using constants from
    riscv_internal_types

    Any output ports driven by these signals are simple wires, of
    course.

    All base instruction types (R/I/S/U) need the opcode @combs.opc
    field; for those that require rd, rs1 and rs2 they is always in
    the same place; the remaining fields are funct3 (used in R/I/S
    types), funct7 (used in R type instructions), and various
    immediate fields.

    Spec 2.2 fig 2.3 shows opcode (must_be_ones and opc); rd, rs1, rs2; funct3 and funct7.
    The other fields in fig 2.3 relate to the immediate value (see immediate_decode)
    """: {
        combs.use_debug = instruction.debug.valid;
        if (rv_cfg_debug_force_disable || !riscv_config.debug_enable) {
            combs.use_debug = 0;
        }

        /*b  Break out the instruction word */
        combs.must_be_ones  = instruction.data[ 2;riscv_i32_ones]; // 2;0
        combs.opc           = instruction.data[ 5;riscv_i32_opc ]; // 5;2 - major opcode, table 19.1
        idecode_inst.rd          = instruction.data[ 5;riscv_i32_rd  ]; // 5;7
        combs.funct3        = instruction.data[ 3;riscv_i32_f3  ]; // 3;12
        idecode_inst.rs1         = instruction.data[ 5;riscv_i32_rs1 ]; // 5;15
        idecode_inst.rs2         = instruction.data[ 5;riscv_i32_rs2 ]; // 5;20
        combs.funct7        = instruction.data[ 7;riscv_i32_f7  ]; //  7;25
    }

    /*b Decode the immediate value
     */
    immediate_decode """
    Decode the immediate value based on the instruction opcode class.

    The immediate is generally a sign-extended value, with the sign
    bit coming from the top bit of the instruction.  Hence @a
    combs.imm_signed is created as a 32 bit value of either all ones
    or all zeros, to be used as a sign extension bit vector as required.

    The immediate variants of the RISC-V I32 base instruction (fig 2.4) are:

      I-type (12-bit sign extended using i[31], i[11;20]) (register-immediate, load, jalr)

      S-type (12-bit sign extended using i[31], i[6;25], i[5;7]) (store)

      B-type ?(13-bit, one zero, sign extended using i[31], i[7], i[6;25], i[4;8], 0) (branch)

      U-type ?(32-bit, twelve zeros, sign extended using i[31]; i[19;12], 12b0 (lui, auipc)

      J-type ?(12-bit sign extended using i[31], i[8;12], i[20], i[10;21], 0) (jal)

    Note that all are sign extended, hence i[31] is replicated on the top bits.
    """: {

        /*b Defaults for the decode */
        combs.imm_signed = combs.funct7[6] ? -1:0;
        idecode_inst.immediate_valid=0;
        idecode_inst.immediate_shift = idecode_inst.rs2;
        idecode_inst.immediate       = bundle(combs.imm_signed[20;0], combs.funct7, idecode_inst.rs2);

        /*b Decode immediate and whether it is used based on instruction class */
        part_switch(combs.opc) {
        case riscv_opc_op_imm, riscv_opc_load, riscv_opc_jalr: { // i format = uses funct7, rs2
            idecode_inst.immediate_valid=1;
        }
        case riscv_opc_store: { // s format - uses funct7, rd (5)
            idecode_inst.immediate_valid=1;
            idecode_inst.immediate = bundle(combs.imm_signed[20;0], combs.funct7, idecode_inst.rd);
        }
        case riscv_opc_branch: { // sb format - uses funct7[6], rd[0], funct7[6;0], rd[4;1], 1b0
            idecode_inst.immediate_valid=1;
            idecode_inst.immediate = bundle(combs.imm_signed[19;0], combs.funct7[6], idecode_inst.rd[0], combs.funct7[6;0], idecode_inst.rd[4;1], 1b0);
        }
        case riscv_opc_jal: { // uj format - uses funct7[6], rs1 (5), funct3 (3), rs2[0], funct7[6;0], rs2[4;1], 1b0
            idecode_inst.immediate_valid=1;
            idecode_inst.immediate = bundle(combs.imm_signed[11;0], combs.funct7[6], idecode_inst.rs1, combs.funct3, idecode_inst.rs2[0], combs.funct7[6;0], idecode_inst.rs2[4;1], 1b0);
        }
        case riscv_opc_lui, riscv_opc_auipc: { // u format - uses funct7, rs2, rs1, funct3, 12b0
            idecode_inst.immediate_valid=1;
            idecode_inst.immediate = bundle(combs.funct7, idecode_inst.rs2, idecode_inst.rs1, combs.funct3, 12b0);
        }
        case riscv_opc_system: {
            idecode_inst.immediate_valid = instruction.data[14]; // for csr write immediates only, data written is rs1
            idecode_inst.immediate       = bundle(27b0, idecode_inst.rs1);
        }
        }
    }

    /*b CSR access decode - debug or not regular */
    csr_access_decode: {
        csr_access = {*=0};
        csr_access.address = instruction.data[12;20];
        csr_access.mode    = instruction.mode;
        csr_access.access  = riscv_csr_access_none;
        part_switch (combs.funct3[2;0]) {
        case riscv_f3_csrrw:      {
            csr_access.access = riscv_csr_access_rw;
            if (idecode_inst.rd==0) { csr_access.access = riscv_csr_access_write; } // True for CSRRW and CSRRWI
        }
        case riscv_f3_csrrs:      {
            csr_access.access = riscv_csr_access_rs;
            if (!combs.rs1_nonzero) { csr_access.access = riscv_csr_access_read; } // True for CSRRS and CSRRSI
        }
        case riscv_f3_csrrc:      {
            csr_access.access = riscv_csr_access_rc;
            if (!combs.rs1_nonzero) { csr_access.access = riscv_csr_access_read; } // True for CSRRC and CSRRCI
        }
        }
        if (combs.use_debug) {
            csr_access.mode    = rv_mode_debug;
            csr_access.address = instruction.debug.data[12;0];
            if (!instruction.debug.data[12]) { // CSRs have bit 12 clear
                csr_access.access  = riscv_csr_access_read;
                if (instruction.debug.debug_op==rv_inst_debug_op_write_reg) {
                    csr_access.access  = riscv_csr_access_write;
                }
            }
        }
        riscv_csrs_decode csrs_decode_i32( csr_access <= csr_access,
                                           csr_decode => csr_decode );
    }

    /*b Basic instruction decode
     */
    instruction_decode """
    Decode the instruction
    """: {
        /*b  Defaults */
        idecode_inst.ext = {*=0};
        idecode_inst.is_compressed = 0;
        idecode_inst.rs1_valid = 0;
        idecode_inst.rs2_valid = 0;
        idecode_inst.rd_written = 0;
        idecode_inst.csr_access = csr_access;
        idecode_inst.csr_access.access = riscv_csr_access_none;
        idecode_inst.csr_access.select = csr_decode.csr_select;

        /*b Decode 'opc' */
        combs.is_imm_op = (combs.opc==riscv_opc_op_imm);
        idecode_inst.op = riscv_op_illegal;
        idecode_inst.illegal = 1;
        idecode_inst.subop = riscv_subop_valid; // so only opc has to be set to 'valid'
        idecode_inst.funct7 = combs.funct7;
        combs.rs1_nonzero = (idecode_inst.rs1 != 0);

        //riscv_shift_op_count               = 4b1010,
        idecode_inst.shift_op = riscv_shift_op_left_logical_zeros;
        full_switch (combs.funct7[2;5]) {
        case 2b00: { idecode_inst.shift_op = (combs.funct3==riscv_f3_sll) ? riscv_shift_op_left_logical_zeros : riscv_shift_op_right_logical_zeros; }
        case 2b01: { idecode_inst.shift_op = (combs.funct3==riscv_f3_sll) ? riscv_shift_op_left_logical_zeros : riscv_shift_op_right_arithmetic;    }
        case 2b10: { idecode_inst.shift_op = (combs.funct3==riscv_f3_sll) ? riscv_shift_op_left_rotate        : riscv_shift_op_right_rotate;        }
        case 2b11: { idecode_inst.shift_op = (combs.funct3==riscv_f3_sll) ? riscv_shift_op_left_logical_ones  : riscv_shift_op_right_logical_ones;  }
        }
        if (rv_cfg_i32_bitmap_enhanced_shift_enable) {
            part_switch (combs.funct7[4;3]) { // 4b0000, 4b0100 standard; 4b0001 muldiv
            case 4b0000: { idecode_inst.shift_op = (combs.funct3==riscv_f3_sll) ? riscv_shift_op_left_logical_zeros : riscv_shift_op_right_logical_zeros;  }
            case 4b0100: { idecode_inst.shift_op = (combs.funct3==riscv_f3_sll) ? riscv_shift_op_left_logical_zeros : riscv_shift_op_right_arithmetic;  }
            case 4b1000: { idecode_inst.shift_op = (combs.funct3==riscv_f3_sll) ? riscv_shift_op_left_logical_ones  : riscv_shift_op_right_logical_ones;  }
            case 4b1001: { idecode_inst.shift_op = (combs.funct3==riscv_f3_sll) ? riscv_shift_op_left_rotate        : riscv_shift_op_right_rotate;  }
            case 4b1010: { idecode_inst.shift_op = (combs.funct3==riscv_f3_sll) ? riscv_shift_op_reverse            : riscv_shift_op_count;  }
            case 4b1100: { idecode_inst.shift_op = (combs.funct3==riscv_f3_sll) ? riscv_shift_op_byte_insert        : riscv_shift_op_byte_insert;  }
            }
        }

        part_switch (combs.opc) {
        case riscv_opc_lui:    { // load upper immediate, uses u format
            // Spec 2.2 section 2.4
            idecode_inst.op = riscv_op_lui;
            idecode_inst.rd_written = 1;
            idecode_inst.illegal = 0;
        }
        case riscv_opc_auipc:  { // add upper immediate pc, uses u format
            // Spec 2.2 section 2.4
            idecode_inst.op = riscv_op_auipc;
            idecode_inst.rd_written = 1;
            idecode_inst.illegal = 0;
        }
        case riscv_opc_jal:    { // jump-and-link, uses uj format
            // Spec 2.2 section 2.5
            // Note that JAL is potentially an unconditional decode-time branch
            idecode_inst.op = riscv_op_jal;
            idecode_inst.rd_written = 1; // Note rd==0 (J rather than JAL) clears this later
            idecode_inst.illegal = 0;
        }
        case riscv_opc_jalr:   { // jump-and-link register, uses i format
            // Spec 2.2 section 2.5
            // Note that JALR is an ALU-time branch
            idecode_inst.op = riscv_op_jalr;
            idecode_inst.rs1_valid = 1;
            idecode_inst.rd_written = 1; // Note rd==0 (J rather than JAL) clears this later
            idecode_inst.illegal = 0;
        }
        case riscv_opc_load:   { // load rd from rs1+offset, uses i format
            // Spec 2.2 section 2.6
            idecode_inst.op = riscv_op_mem;
            idecode_inst.subop = bundle(1b0, combs.funct3);
            idecode_inst.rs1_valid = 1;
            idecode_inst.rd_written = 1;
            idecode_inst.illegal = 0;
        }
        case riscv_opc_store:  { // store rs2 at rs1+offset, uses s format
            // Spec 2.2 section 2.6
            idecode_inst.op = riscv_op_mem;
            idecode_inst.subop = bundle(1b1, combs.funct3);
            idecode_inst.rs1_valid = 1;
            idecode_inst.rs2_valid = 1;
            idecode_inst.illegal = 0;
        }
        case riscv_opc_branch: { // branch if rs1 <=> rs2 to pc+imm, uses sb format, conditional branch to +-4kB
            // Spec 2.2 section 2.5
            // Note that Bxx is an ALU-time branch
            idecode_inst.op = riscv_op_branch;
            idecode_inst.rs1_valid = 1;
            idecode_inst.rs2_valid = 1;
            idecode_inst.subop = riscv_subop_illegal;
            idecode_inst.illegal = 0;
            part_switch (combs.funct3) {
            case riscv_f3_beq:  { idecode_inst.subop = riscv_subop_beq;  }
            case riscv_f3_bne:  { idecode_inst.subop = riscv_subop_bne;  }
            case riscv_f3_blt:  { idecode_inst.subop = riscv_subop_blt;  }
            case riscv_f3_bltu: { idecode_inst.subop = riscv_subop_bltu; }
            case riscv_f3_bge:  { idecode_inst.subop = riscv_subop_bge;  }
            case riscv_f3_bgeu: { idecode_inst.subop = riscv_subop_bgeu; }
            }
        }
        case riscv_opc_op, riscv_opc_op_imm: { // rd = rs1 op rs2/imm, uses r or i format
            // Spec 2.2 section 2.4
            idecode_inst.op = riscv_op_alu;
            idecode_inst.rs1_valid = 1;
            idecode_inst.rs2_valid = !combs.is_imm_op;
            idecode_inst.rd_written = 1;
            if ((combs.funct7==1) && (!combs.is_imm_op)){
                if ((rv_cfg_i32m_force_disable==0) && riscv_config.i32m) {
                    idecode_inst.illegal = 0;
                    idecode_inst.op = riscv_op_muldiv;
                    full_switch (combs.funct3) {
                    case riscv_f3_mul:    { idecode_inst.subop = riscv_subop_mull; }
                    case riscv_f3_mulh:   { idecode_inst.subop = riscv_subop_mulhss; }
                    case riscv_f3_mulhsu: { idecode_inst.subop = riscv_subop_mulhsu; }
                    case riscv_f3_mulhu:  { idecode_inst.subop = riscv_subop_mulhu; }
                    case riscv_f3_div:    { idecode_inst.subop = riscv_subop_divs; }
                    case riscv_f3_divu:   { idecode_inst.subop = riscv_subop_divu; }
                    case riscv_f3_rem:    { idecode_inst.subop = riscv_subop_rems; }
                    case riscv_f3_remu:   { idecode_inst.subop = riscv_subop_remu; }
                    }
                }
            } else {
                idecode_inst.illegal = (!combs.is_imm_op) && (combs.funct7!=0) && (combs.funct7!=0x20);
                full_switch (combs.funct3) {
                case riscv_f3_addsub: { idecode_inst.subop = (!combs.is_imm_op && combs.funct7[5]) ? riscv_subop_sub : riscv_subop_add; }
                case riscv_f3_slt:    { idecode_inst.subop = riscv_subop_slt; }
                case riscv_f3_sltu:   { idecode_inst.subop = riscv_subop_sltu; }
                case riscv_f3_xor :   { idecode_inst.subop = riscv_subop_xor; }
                case riscv_f3_or:     { idecode_inst.subop = riscv_subop_or; }
                case riscv_f3_and:    { idecode_inst.subop = riscv_subop_and; }
                case riscv_f3_sll:    {
                    idecode_inst.illegal = (combs.funct7!=0);
                    idecode_inst.subop   = riscv_subop_sll;
                    if (rv_cfg_i32_bitmap_enhanced_shift_enable) {
                        if (combs.funct7[6]) { idecode_inst.illegal = 0; } // bit manip extension legalizes all f7[6] set
                    }
                }
                case riscv_f3_srlsra: {
                    idecode_inst.illegal = ((combs.funct7!=0) &&(combs.funct7!=7b0100000));
                    idecode_inst.subop   =  riscv_subop_srla; // SRAI has funct7[5] set, else SRLI
                    if (rv_cfg_i32_bitmap_enhanced_shift_enable) {
                        if (combs.funct7[6]) { idecode_inst.illegal = 0; } // bit manip extension legalizes all f7[6] set
                    }
                }
                default:          {
                    idecode_inst.illegal = 1;
                }
                }
            }
        }
        case riscv_opc_misc_mem: { // uses i format
            // Spec 2.2 section 2.7
            idecode_inst.illegal = 0;
            idecode_inst.op = riscv_op_misc_mem;
            idecode_inst.subop = combs.funct3[0] ? riscv_subop_fence_i : riscv_subop_fence;
        }
        case riscv_opc_system: { // system access, or csr rw/rs/rc - uses i format
            // Spec 2.2 section 2.8
            idecode_inst.op = riscv_op_system;
            idecode_inst.rs1_valid = 1;
            idecode_inst.rd_written = 1;
            idecode_inst.csr_access.access = csr_access.access;
            idecode_inst.illegal           = csr_decode.illegal_access; // valid based on access which is okay for non-CSR instructions
            full_switch (combs.funct3[2;0]) {
            case riscv_f3_csrrw: { idecode_inst.op = riscv_op_csr; idecode_inst.subop = riscv_subop_csrrw; }
            case riscv_f3_csrrs: { idecode_inst.op = riscv_op_csr; idecode_inst.subop = riscv_subop_csrrs; }
            case riscv_f3_csrrc: { idecode_inst.op = riscv_op_csr; idecode_inst.subop = riscv_subop_csrrc; }
            case riscv_f3_privileged: {
                idecode_inst.op = riscv_op_system;
                full_switch (instruction.data[12;20]) {
                case riscv_f12_ecall:  { idecode_inst.subop = riscv_subop_ecall;  }
                case riscv_f12_ebreak: { idecode_inst.subop = riscv_subop_ebreak; }
                case riscv_f12_mret:   {
                    idecode_inst.subop = riscv_subop_mret;
                    idecode_inst.illegal = (instruction.mode < rv_mode_machine);
                }
                case riscv_f12_mwfi:   {
                    idecode_inst.subop = riscv_subop_mwfi;
                    idecode_inst.illegal = (instruction.mode < rv_mode_machine);
                }
                default:  { idecode_inst.illegal = 1; }
                }
            }
            }
        }
        case riscv_opc_custom_0: {
            if (rv_cfg_i32_custom0_enable==1) {
                idecode_inst.illegal = 0;
                idecode_inst.op = riscv_op_custom_0;
                idecode_inst.subop = bundle(1b0,combs.funct3);
                idecode_inst.rs1_valid = 1;
                if (rv_cfg_i32_custom0_as_load==1)  {idecode_inst.rs2_valid = 1;}
                if (rv_cfg_i32_custom0_as_store==1) {idecode_inst.rd_written = 1;}
            }
        }
        case riscv_opc_custom_1: {
            if (rv_cfg_i32_custom1_enable==1) {
                idecode_inst.illegal = 0;
                idecode_inst.op = riscv_op_custom_1;
                idecode_inst.subop = bundle(1b0,combs.funct3);
                idecode_inst.rs1_valid = 1;
                if (rv_cfg_i32_custom1_as_load==1)  {idecode_inst.rs2_valid = 1;}
                if (rv_cfg_i32_custom1_as_store==1) {idecode_inst.rd_written = 1;}
            }
        }
        case riscv_opc_custom_2: {
            if (rv_cfg_i32_custom2_enable==1) {
                idecode_inst.illegal = 0;
                idecode_inst.op = riscv_op_custom_2;
                idecode_inst.subop = bundle(1b0,combs.funct3);
                idecode_inst.rs1_valid = 1;
                if (rv_cfg_i32_custom2_as_load==1)  {idecode_inst.rs2_valid = 1;}
                if (rv_cfg_i32_custom2_as_store==1) {idecode_inst.rd_written = 1;}
            }
        }
        case riscv_opc_custom_3: {
            if (rv_cfg_i32_custom3_enable==1) {
                idecode_inst.illegal = 0;
                idecode_inst.op = riscv_op_custom_3;
                idecode_inst.subop = bundle(1b0,combs.funct3);
                idecode_inst.rs1_valid = 1;
                if (rv_cfg_i32_custom3_as_load==1)  {idecode_inst.rs2_valid = 1;}
                if (rv_cfg_i32_custom3_as_store==1) {idecode_inst.rd_written = 1;}
            }
        }
        }

        if (combs.must_be_ones != -1) { // rv32i 32-bit encodings only
            idecode_inst.illegal = 1;
        }
        if (idecode_inst.rs1 == 0) {
            idecode_inst.rs1_valid = 0;
        }
        if (idecode_inst.rs2 == 0) {
            idecode_inst.rs2_valid = 0;
        }
        if (idecode_inst.rd == 0) {
            idecode_inst.rd_written = 0;
        }

        if (riscv_config.e32 || rv_cfg_e32_force_enable) {
            if (idecode_inst.rs1_valid && idecode_inst.rs1[4]) {
                idecode_inst.illegal = 1;
            }
            if (idecode_inst.rs2_valid && idecode_inst.rs2[4]) {
                idecode_inst.illegal = 1;
            }
            if (idecode_inst.rd_written && idecode_inst.rd[4]) {
                idecode_inst.illegal = 1;
            }
        }
    }

    /*b Debug instruction decode */
    debug_decode : {
        idecode_debug = {*=0};
        idecode_debug.immediate = instruction.data;
        idecode_debug.rs1       = instruction.debug.data[5;0];
        idecode_debug.rs1_valid = 1;
        idecode_debug.rs2       = 0;
        idecode_debug.rs2_valid = 0;
        idecode_debug.rd        = instruction.debug.data[5;0];
        idecode_debug.rd_written = 0;
        idecode_debug.immediate_valid = 1;
        idecode_debug.op    = riscv_op_alu;
        idecode_debug.subop = riscv_subop_or; // alu_result = rs1 | rs2_or_imm
        idecode_debug.csr_access.access  = riscv_csr_access_none;
        idecode_debug.csr_access.address = instruction.debug.data[12;0];
        idecode_debug.csr_access.select  = csr_decode.csr_select;
        if (instruction.debug.data[12]) { // GPR access
            full_switch (instruction.debug.debug_op) {
            case rv_inst_debug_op_read_reg: {
                idecode_debug.rs1_valid       = 0;
                idecode_debug.immediate_valid = 0;
            }
            case rv_inst_debug_op_write_reg: { // rd <= 0 | imm
                idecode_debug.rs1             = 0;
                idecode_debug.rs1_valid       = 0;
                idecode_debug.immediate_valid = 1;
                idecode_debug.rd_written      = 1;
            }
            }
        } else { // CSR access
            idecode_debug.op    = riscv_op_csr;
            idecode_debug.subop = riscv_subop_or; // csr read
            full_switch (instruction.debug.debug_op) {
            case rv_inst_debug_op_read_reg: {
                idecode_debug.csr_access.access = riscv_csr_access_read;
                idecode_debug.rs1_valid       = 0;
                idecode_debug.immediate_valid = 0;
            }
            case rv_inst_debug_op_write_reg: { // csr write
                idecode_debug.csr_access.access = riscv_csr_access_write;
                idecode_debug.rs1_valid       = 0;
                idecode_debug.immediate_valid = 1;
            }
            }
        }
    }

    /*b Select output from debug or regular */
    select_output : {
        idecode = idecode_inst;
        if (combs.use_debug) {
            idecode = idecode_debug;
        }
    }

    /*b All done */
}
