/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   riscv_minimal.cdl
 * @brief  Minimal RISC-V implementation ported to CDL
 *
 * CDL implementation of minimal RISC-V teaching implementation
 *
 * This is a two-stage pipeline implementation, with instruction fetch
 * of the next PC occuring simultaneously with the decode, register
 * read, ALU, data read/write request, data read memory access, and
 * register update.
 *
 * The instruction memory request, then, becomes valid dependent on
 * the decode of the registered instruction last fetched. For most
 * branches this requires only a small amount of logic, but for
 * jump-and-link-register instructions (which uses the full ALU
 * result) this may take a considerable amount of gates to determine
 * the correct branch target and hence next instruction fetch.  Hence
 * the instruction memory request is valid after a considerable delay
 * from the start of the cycle.
 *
 * The return value from the instruction memory request must be valid
 * before the end of the cycle.
 *
 * Any instruction memory implementation must start its access well
 * after the CPU clock edge, , as the request is valid after the CPU
 * clock edge; the resultant read data delay (from the clock edge)
 * then has to be factored in to determine when the next CPU clock
 * edge can occur. Hence it may be sensible to use a double speed
 * clock (e.g. 'fast_clk') to generate CPU clock edges (every other
 * fast_clk edge) and SRAM access clock edges (for a synchronous
 * memory) on the intervening fast_clk edges.
 *
 * The data memory request becomes valid, again, a fair time after the
 * CPU clock edge, as it requires instruction decode, register fetch,
 * and ALU operation to occur prior to the memory address being valid.
 *
 * The data memory response must be valid (for read data!) in the same
 * CPU cycle, as the returning data has to be rotated to the correct
 * byte lanes and prepared for the register file write.
 *
 * Hence a data memory implementation can be similar to that proposed
 * for the instruction memory - that is, accesses start on a memory
 * clock edge that is in the middle of a CPU clock edge, by using a
 * fast_clk.
 *
 */

/*a Includes
 */
include "cpu/riscv/riscv.h"
include "cpu/riscv/riscv_modules.h"

/*a Module
 */
module riscv_minimal_debug( clock clk,
                            input bit reset_n,
                            output t_riscv_mem_access_req  dmem_access_req,
                            input  t_riscv_mem_access_resp dmem_access_resp,
                            output t_riscv_fetch_req       ifetch_req,
                            input  t_riscv_fetch_resp      ifetch_resp,
                            input  t_riscv_debug_mst       debug_mst "Driven by debug module to all RISC-V cores",
                            output t_riscv_debug_tgt       debug_tgt "Wired-or response bus from all RISC-V cores",

                            input  t_riscv_config          riscv_config,
                            input bit[6] rv_select,
                            output t_riscv_i32_trace       trace
)
"""
"""
{

    /*b State and comb
     */
    net t_riscv_fetch_req       pipeline_ifetch_req;
    net t_riscv_fetch_resp      pipeline_ifetch_resp;
    net t_riscv_fetch_req       ifetch_req;
    net t_riscv_mem_access_req  dmem_access_req;
    net t_riscv_i32_coproc_controls  coproc_controls;
    comb t_riscv_i32_coproc_response   coproc_response;
    net t_riscv_i32_trace       trace;
    net t_riscv_pipeline_debug_control debug_control;
    net t_riscv_pipeline_debug_response debug_response;
    net t_riscv_debug_tgt       debug_tgt;

    /*b Pipeline and debug */
    pipeline_debug: {
        coproc_response = {*=0};
        riscv_i32_ifetch_debug  ifetch_debug( pipeline_ifetch_req <= pipeline_ifetch_req,
                                              pipeline_ifetch_resp => pipeline_ifetch_resp,
                                              pipeline_trace <= trace,
                                              debug_control <= debug_control,
                                              debug_response => debug_response,
                                              ifetch_req => ifetch_req,
                                              ifetch_resp <= ifetch_resp );

        riscv_i32_pipeline_debug pdm( clk <- clk,
                                      reset_n <= reset_n,
                                      debug_mst <= debug_mst,
                                      debug_tgt => debug_tgt,
                                      debug_control => debug_control,
                                      debug_response <= debug_response,
                                      rv_select <= rv_select );

        // Pipeline must contain CSRs that include the debug CSRs (riscv_config must enable debug?)
        riscv_i32c_pipeline pipeline(clk <- clk,
                                     reset_n <= reset_n,
                                     ifetch_req => pipeline_ifetch_req,
                                     ifetch_resp <= pipeline_ifetch_resp,
                                     dmem_access_req => dmem_access_req,
                                     dmem_access_resp <= dmem_access_resp,
                                     coproc_controls => coproc_controls,
                                     coproc_response <= coproc_response,
                                     riscv_config <= riscv_config,
                                     trace => trace );
    }

    /*b All done */
}

