/** Copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *   http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * @file   bbc_micro_with_rams.cdl
 * @brief  BBC microcomputer with RAMs module
 *
 * CDL implementation of a BBC microcomputer with RAMs for framebuffer
 * and display; this is suitable for instantiation in an FPGA.
 *
 */
/*a Includes */
include "microcomputers/bbc/bbc_types.h"
include "microcomputers/bbc/bbc_submodules.h"
include "video/framebuffer_modules.h"
include "srams.h"

/*a Module */
module bbc_micro_with_rams( clock clk "4MHz clock in as a minimum",
                            clock video_clk,
                            input bit reset_n,
                            input t_csr_request csr_request,
                            output t_csr_response csr_response,
                            input t_bbc_micro_sram_request   host_sram_request,
                            output t_bbc_micro_sram_response host_sram_response,
                            output t_bbc_display_sram_write display_sram_write,
                            output t_video_bus video_bus )
{
    net t_video_bus video_bus;
    net t_bbc_display display;
    net  bit keyboard_reset_n;
    net t_bbc_floppy_op floppy_op;
    net  t_bbc_floppy_response floppy_response;

    net t_bbc_clock_status clock_status;
    net t_bbc_clock_control clock_control;
    net t_csr_response clocking_csr_response;
    net t_csr_response display_sram_csr_response;
    net t_csr_response keyboard_csr_response;
    net t_csr_response floppy_sram_csr_response;
    net t_csr_response framebuffer_csr_response;

    net t_bbc_floppy_sram_request floppy_sram_request;
    net t_bbc_floppy_sram_response floppy_sram_response;
    net t_bbc_display_sram_write display_sram_write;

    net t_bbc_micro_sram_request bbc_micro_host_sram_request;
    net t_bbc_micro_sram_response bbc_micro_host_sram_response;
    net t_bbc_micro_sram_response host_sram_response;
    
    gated_clock clock clk active_high enable_clk_2MHz_video   clk_2MHz_video_clock "Clock that mirrors 2MHz falling -  video data from RAM is valid at this edge, so used by CRTC, SAA5050 latches, SAA5050, vidproc";
    gated_clock clock clk active_high enable_cpu_clk          clk_cpu  "6502 clock, >=2MHz but extended when accessing 1MHz peripherals";
    comb bit enable_clk_2MHz_video;
    comb bit enable_cpu_clk;

    // FDC clocks off rising CPU clock
    // display clocks off falling 2MHz clock
    //
    comb bit bbc_reset_n;
    net t_bbc_keyboard keyboard;
    comb t_sram_access_req display_sram_access_req;
    stuff """
    """: {
        csr_response = floppy_sram_csr_response;
        csr_response |= display_sram_csr_response;
        csr_response |= clocking_csr_response;
        csr_response |= keyboard_csr_response;
        enable_clk_2MHz_video   = clock_control.enable_2MHz_video; // used for clock enable and to choose which source of SRAM read
        enable_cpu_clk          = clock_control.enable_cpu;
        bbc_micro_clocking clocking( clk <- clk,
                                     reset_n <= reset_n,
                                     clock_status <= clock_status,
                                     clock_control => clock_control,
                                     csr_request <= csr_request,
                                     csr_response => clocking_csr_response );

        bbc_reset_n = reset_n & !clock_control.reset_cpu;
        bbc_micro bbc(clk <- clk,
                      reset_n <= bbc_reset_n,
                      clock_control <= clock_control,
                      clock_status  => clock_status,
                      keyboard <= keyboard,
                      display => display,
                      keyboard_reset_n => keyboard_reset_n,
                      floppy_op => floppy_op,
                      floppy_response <= floppy_response,
                      host_sram_request <= bbc_micro_host_sram_request,
                      host_sram_response => bbc_micro_host_sram_response
            );
    
        bbc_display_sram display_sram( clk <- clk_2MHz_video_clock,
                                       reset_n <= reset_n,
                                       display <= display,
                                       sram_write => display_sram_write,
                                       csr_request <= csr_request,
                                       csr_response => display_sram_csr_response
            );

        bbc_keyboard_csr keyboard_csr( clk <- clk_cpu,
                                       reset_n <= reset_n,
                                       keyboard => keyboard,
                                       keyboard_reset_n <= 1b1, // not really used in this model - comes from CSRs
                                       csr_request <= csr_request,
                                       csr_response => keyboard_csr_response
            );

        bbc_floppy_sram floppy_sram( clk <- clk_cpu, // FDC interacts with floppy at cpu clock
                                     reset_n <= reset_n,
                                     floppy_op <= floppy_op,
                                     csr_request <= csr_request,
                                     floppy_response => floppy_response,
                                     sram_request => floppy_sram_request,
                                     sram_response <= floppy_sram_response,
                                     csr_response => floppy_sram_csr_response
            );

        bbc_micro_rams rams( clk <- clk,
                             reset_n <= reset_n,
                             clock_control <= clock_control,
                             host_sram_request <= host_sram_request,
                             host_sram_response => host_sram_response,
                             display_sram_write <= display_sram_write,
                             floppy_sram_request <= floppy_sram_request,
                             floppy_sram_response => floppy_sram_response,
                             bbc_micro_host_sram_request => bbc_micro_host_sram_request,
                             bbc_micro_host_sram_response <= bbc_micro_host_sram_response );

        display_sram_access_req = {*=0};
        display_sram_access_req.valid      = display_sram_write.enable;
        display_sram_access_req.address    = bundle(16b0,display_sram_write.address);
        display_sram_access_req.write_data = bundle(16b0,display_sram_write.data);
        framebuffer fb( csr_clk <- clk_cpu,
                        sram_clk <- clk_2MHz_video_clock,
                        video_clk <- video_clk,
                        reset_n <= reset_n,
                        video_bus => video_bus,
                        display_sram_write <= display_sram_access_req,
                        csr_request <= csr_request,
                        csr_response => framebuffer_csr_response
            );
                        
    }
}
