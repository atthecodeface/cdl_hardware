/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   riscv_i32_decode.cdl
 * @brief  Instruction decoder for RISC-V implementation
 *
 * CDL implementation of RISC-V instruction decode based on the RISC-V
 * specification v2.1.
 *
 */

/*a Includes
 */
include "riscv_internal_types.h"
include "riscv_submodules.h"
include "riscv.h"

/*a Module
 */
module riscv_e32c_decode( input t_riscv_i32_inst    instruction,
                          output t_riscv_i32_decode idecode,
                          input  t_riscv_config     riscv_config
)
"""
Instruction decoder for RISC-V RV32E instruction set.

This is based on the RISC-V v2.1 specification (hence figure numbers
are from that specification)
"""
{
    net t_riscv_i32_decode rv32i_idecode;

    /*b Basic instruction decode - RV32I
     */
    instruction_decode """
    Decode the instruction
    """: {
        riscv_i32c_decode rv32ic_decode( instruction <= instruction,
                                       idecode => rv32i_idecode,
                                       riscv_config <= riscv_config );

        idecode = rv32i_idecode;
        if (rv32i_idecode.rs1_valid && rv32i_idecode.rs1[4]) {
            idecode.illegal = 1;
        }
        if (rv32i_idecode.rs2_valid && rv32i_idecode.rs2[4]) {
            idecode.illegal = 1;
        }
        if (rv32i_idecode.rd_written && rv32i_idecode.rd[4]) {
            idecode.illegal = 1;
        }

        /*b All done */
    }

    /*b All done */
}
