/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   tb_riscv_minimal.cdl
 * @brief  Testbench for minimal RISC-V
 *
 */

/*a Includes
 */
include "srams.h"
include "types/apb.h"
include "apb/apb_targets.h"
include "cpu/riscv/riscv.h"
include "cpu/riscv/riscv_modules.h"
include "cpu/riscv/riscv_pipeline.h"
include "cpu/riscv/riscv_submodules.h"
include "cpu/riscv/chk_riscv.h"

/*a Types */
/*t t_drop_data */
typedef enum[2] {
    drop_data_none,
    drop_data_16,
    drop_data_32,
    drop_data_all
} t_drop_data;

/*t t_sram_request */
typedef struct {
    bit     valid;
    bit     read_not_write;
    bit[32] address;
    bit[4]  byte_enable;
    bit[32] write_data;
} t_sram_request;

/*t t_inst_combs */
typedef struct {
    bit[64] data_before_drop;
    bit[64] data_after_drop;
    bit[4] half_words_valid;
    bit[4] half_words_will_be_valid;
    t_sram_request sram_request;
    bit request_initial_half;
    t_drop_data drop_data;
} t_inst_combs;

/*t t_inst_state */
typedef struct {
    bit[4]  half_words_valid_before_reading;
    bit     sram_reading;
    bit     initial_half;
    bit[32] address;
    bit[64] data;
} t_inst_state;

/*t t_data_combs */
typedef struct {
    t_sram_request sram_request;
    bit apb_request_valid;
} t_data_combs;

/*t t_data_state */
typedef struct {
    t_riscv_mem_access_req dmem_access_in_progress;
    t_apb_request apb;
} t_data_state;

/*t t_arbiter_combs */
typedef struct {
    t_sram_request sram_request;
    bit grant_to_inst;
    bit grant_to_data;
} t_arbiter_combs;

/*a External modules */
extern module se_test_harness( clock clk, output t_jtag jtag, output bit tck_enable, input bit tdo )
{
    timing from rising clock clk jtag, tck_enable;
    timing to rising clock clk tdo;
}

/*a Module
 */
module tb_riscv_i32mc_system( clock jtag_tck,
                                 clock clk,
                                 input bit reset_n
)
{
    /*b Default clock and reset
     */
    default clock clk;
    default reset active_low reset_n;

    /*b Configuration and tie-offs
     */
    clocked t_riscv_config riscv_config={*=0, i32c=1, i32m=1, i32m_fuse=1, coproc_disable=0, debug_enable=1} ;
    clocked t_riscv_irqs                 irqs= {*=0};
    clocked t_timer_control timer_control = {*=0};

    /*b Nets
     */
    net t_jtag jtag;
    net bit tdo;
    net bit[5]ir;
    net t_jtag_action dr_action;
    net bit[50]dr_in;
    net bit[50]dr_tdi_mask;
    net bit[50]dr_out;
    net bit tck_enable;
    comb bit tck_enable_fix;
    gated_clock clock jtag_tck active_high tck_enable_fix jtag_tck_gated;

    net   t_apb_request  dm_apb_request  "APB request for debug";
    net   t_apb_response dm_apb_response "APB response for debug";
    net   t_riscv_debug_mst debug_mst;
    comb  t_riscv_debug_tgt debug_tgt;
    net   t_riscv_debug_tgt debug_tgt0;

    net  t_riscv_mem_access_req  dmem_access_req;
    comb t_riscv_mem_access_resp dmem_access_resp;

    net  t_riscv_fetch_req  rv_imem_access_req;
    comb t_riscv_fetch_resp rv_imem_access_resp;
    net t_riscv_csr_controls      csr_controls;
    net t_riscv_csr_data          csr_data;
    net t_riscv_csr_access        csr_access;
    net t_riscv_csrs_minimal csrs;

    /*b Nets for the pipeline
     */
    net t_riscv_pipeline_state        pipeline_state;
    net t_riscv_pipeline_control      pipeline_control;
    net t_riscv_pipeline_response     pipeline_response;
    net t_riscv_pipeline_fetch_req    pipeline_fetch_req;
    net t_riscv_pipeline_fetch_data   pipeline_fetch_data;
    net t_riscv_pipeline_trap_request pipeline_trap_request;

    /*b State and comb
     */
    comb    t_inst_combs inst_combs;
    clocked t_inst_state inst_state = {*=0};
    comb    t_data_combs data_combs;
    clocked t_data_state data_state = {*=0};
    comb    t_arbiter_combs arbiter_combs;
    comb    t_apb_request   rv_apb_request;
    comb    t_apb_response  rv_apb_response;
    comb    t_apb_request   timer_apb_request;
    net     t_apb_response  timer_apb_response;
    net     t_timer_value   timer_value;
    net bit[32] sram_read_data;

    net t_riscv_i32_coproc_controls  coproc_controls;
    net t_riscv_i32_coproc_response  coproc_response;
    net t_riscv_i32_coproc_response  pipeline_coproc_response;

    net t_riscv_i32_trace trace;
    comb t_riscv_packed_trace_control trace_control;
    net t_riscv_i32_packed_trace packed_trace;
    net t_riscv_i32_compressed_trace compressed_trace;
    net t_riscv_i32_decompressed_trace decompressed_trace;
    net bit[5] nybbles_consumed;

    /*b Configuration
     */
    configuration """
    Tie-offs are best done as clocked signals, with the reset value and the assigned values being equal.
    In synthesis the flops will be optimized out as tied-low or tied-high.
    """ : {
        riscv_config <= {*=0};
        riscv_config.i32c <= 1;
        riscv_config.e32  <= 0;
        riscv_config.i32m <= 1;
        riscv_config.i32m_fuse <= 1;
        riscv_config.coproc_disable <= 0;
        riscv_config.debug_enable <= 1;

        timer_control <= {*=0};
        timer_control.enable_counter   <= 1;
        timer_control.fractional_adder <= 2;
        timer_control.integer_adder    <= 0;
        irqs <= {*=0};
        irqs.mtip <= timer_value.irq;
    }

    /*b SRAM and arbiter */
    sram_and_arbiter: {
        arbiter_combs.grant_to_inst = 0;
        arbiter_combs.grant_to_data = 0;

        arbiter_combs.sram_request = data_combs.sram_request;
        if (data_combs.sram_request.valid) {
            arbiter_combs.grant_to_data = 1;
            arbiter_combs.sram_request  = data_combs.sram_request;
        } elsif (inst_combs.sram_request.valid) {
            arbiter_combs.grant_to_inst = 1;
            arbiter_combs.sram_request = inst_combs.sram_request;
        } else {
            arbiter_combs.sram_request.valid = 0;
        }
        
        /*b SRAM instance */
        se_sram_srw_16384x32_we8 mem(sram_clock     <- clk,
                                     select         <= arbiter_combs.sram_request.valid,
                                     read_not_write <= arbiter_combs.sram_request.read_not_write,
                                     write_enable   <= arbiter_combs.sram_request.byte_enable,
                                     address        <= arbiter_combs.sram_request.address[14;2],
                                     write_data     <= arbiter_combs.sram_request.write_data,
                                     data_out       => sram_read_data );
    }

    /*b Instruction memory
     */
    comb bit riscv_clk_enable;
    srams: {
        riscv_clk_enable = 1;
        /*b Create data buffer value from SRAM read data and current valid data buffer */
        inst_combs.data_before_drop = inst_state.data;
        inst_combs.half_words_valid = inst_state.half_words_valid_before_reading;
        if (inst_state.sram_reading) {
            inst_combs.half_words_valid = inst_state.half_words_valid_before_reading + 2;
            if    (inst_state.half_words_valid_before_reading==0) { inst_combs.data_before_drop[32;0]  = sram_read_data; }
            elsif (inst_state.half_words_valid_before_reading==1) { inst_combs.data_before_drop[32;16] = sram_read_data; }
            else                                                  { inst_combs.data_before_drop[32;32] = sram_read_data; }
            assert (inst_state.half_words_valid_before_reading<=2, "Incorrect value for half_words_valid_before_reading if we are reading");
            if (inst_state.initial_half) {
                inst_combs.data_before_drop[16;0] = sram_read_data[16;16];
                inst_combs.half_words_valid = 1;
            }
        }

        /*b Decode amount of data to drop given request */
        inst_combs.drop_data = drop_data_none;
        full_switch (rv_imem_access_req.req_type) {
        case rv_fetch_none: {
            inst_combs.drop_data = drop_data_all;
        }
        case rv_fetch_nonsequential: {
            inst_combs.drop_data = drop_data_all;
        }
        case rv_fetch_repeat: {
            inst_combs.drop_data = drop_data_none;
        }
        case rv_fetch_sequential_16: {
            inst_combs.drop_data = drop_data_16;
        }
        case rv_fetch_sequential_32: {
            inst_combs.drop_data = drop_data_32;
        }
        }

        /*b Decode amount of data valid after drop */
        inst_combs.half_words_will_be_valid = inst_combs.half_words_valid;
        inst_combs.data_after_drop          = inst_combs.data_before_drop;
        full_switch (inst_combs.drop_data) {
        case drop_data_none: {
            inst_combs.half_words_will_be_valid = inst_combs.half_words_valid;
        }
        case drop_data_16: {
            inst_combs.data_after_drop[48;0] = inst_combs.data_before_drop[48;16];
            if    (inst_combs.half_words_valid==0) { inst_combs.half_words_will_be_valid = 0; }
            elsif (inst_combs.half_words_valid==1) { inst_combs.half_words_will_be_valid = 0; }
            elsif (inst_combs.half_words_valid==2) { inst_combs.half_words_will_be_valid = 1; }
            elsif (inst_combs.half_words_valid==3) { inst_combs.half_words_will_be_valid = 2; }
            else                                   { inst_combs.half_words_will_be_valid = 3; }
        }
        case drop_data_32: {
            inst_combs.data_after_drop[32;0] = inst_combs.data_before_drop[32;32];
            if    (inst_combs.half_words_valid==0) { inst_combs.half_words_will_be_valid = 0; }
            elsif (inst_combs.half_words_valid==1) { inst_combs.half_words_will_be_valid = 0; }
            elsif (inst_combs.half_words_valid==2) { inst_combs.half_words_will_be_valid = 0; }
            elsif (inst_combs.half_words_valid==3) { inst_combs.half_words_will_be_valid = 1; }
            else                                   { inst_combs.half_words_will_be_valid = 2; }
        }
        case drop_data_all: {
            inst_combs.half_words_will_be_valid = 0;
        }
        }

        /*b Decode address to fetch and whether it is valid */
        inst_combs.sram_request = {*=0};
        inst_combs.request_initial_half = 0;
        inst_combs.sram_request.read_not_write  = 1;
        inst_combs.sram_request.address         = inst_state.address;
        full_switch (rv_imem_access_req.req_type) {
        case rv_fetch_none: {
            inst_combs.sram_request.valid = 0;
            inst_combs.request_initial_half  = 0;
        }
        case rv_fetch_nonsequential: {
            inst_combs.sram_request.valid        = 1;
            inst_combs.request_initial_half      = rv_imem_access_req.address[1];
            inst_combs.sram_request.address      = rv_imem_access_req.address;
        }
        default: {
            inst_combs.request_initial_half   = inst_state.initial_half;
            inst_combs.sram_request.valid     = (inst_combs.half_words_will_be_valid<=2);
            inst_combs.sram_request.address   = inst_state.address;
            if (inst_state.sram_reading) {
                inst_combs.request_initial_half   = 0;
                inst_combs.sram_request.address   = inst_state.address+4;
            }
        }
        }

        /*b Present response */
        rv_imem_access_resp          = {*=0};
        rv_imem_access_resp.data     = inst_combs.data_after_drop[32;0];
        if (rv_imem_access_req.req_type!=rv_fetch_none) {
            if (inst_combs.half_words_will_be_valid>=2) {
                rv_imem_access_resp.valid = 1;
            }
        }

        /*b Update state */
        inst_state.data                            <= inst_combs.data_after_drop;
        inst_state.sram_reading                    <= arbiter_combs.grant_to_inst && inst_combs.sram_request.valid;
        inst_state.initial_half                    <= inst_combs.request_initial_half;
        inst_state.half_words_valid_before_reading <= inst_combs.half_words_will_be_valid;
        inst_state.address                         <= inst_combs.sram_request.address;

    }

    /*b Data memory
     */
    data_memory: {
        /*b Decode data request */
        data_combs.apb_request_valid       = 0;
        data_combs.sram_request.valid      = 0;
        data_combs.sram_request.read_not_write = (dmem_access_req.req_type != rv_mem_access_write);
        data_combs.sram_request.address        = dmem_access_req.address;
        data_combs.sram_request.byte_enable    = dmem_access_req.byte_enable;
        data_combs.sram_request.write_data     = dmem_access_req.write_data;
        if (dmem_access_req.valid) {
            data_combs.sram_request.valid          = 1;
            if (dmem_access_req.address[4;28]!=0) { // 3h0xxxxxxx is SRAM, rest is APB
                data_combs.sram_request.valid      = 0;
                data_combs.apb_request_valid       = 1;
            }
        }

        /*b Generate dmem_access_resp and update APB transaction state */
        dmem_access_resp = {*=0};
        dmem_access_resp.ack             = 1;
        dmem_access_resp.access_complete = 1;
        dmem_access_resp.may_still_abort = 0;
        dmem_access_resp.abort_req       = 0;
        dmem_access_resp.read_data       = sram_read_data;
        if (data_state.apb.penable) {
            dmem_access_resp.read_data   = rv_apb_response.prdata;
        }

        if (data_state.apb.psel) {
            dmem_access_resp.ack             = 0;
            dmem_access_resp.access_complete = 0;
            dmem_access_resp.may_still_abort = 1;
            data_state.apb.penable <= 1;
            if (data_state.apb.penable) {
                dmem_access_resp.abort_req = rv_apb_response.perr;
                if (rv_apb_response.pready || rv_apb_response.perr) {
                    dmem_access_resp.ack             = 1;
                    dmem_access_resp.access_complete = 1;
                }
            }
        }

        /*b Update state */
        data_state.dmem_access_in_progress.valid <= 0;
        if (dmem_access_resp.ack) {
            data_state.apb.psel    <= 0;
            data_state.apb.penable <= 0;
            if (dmem_access_req.valid) {
                data_state.dmem_access_in_progress <= dmem_access_req;
                if (data_combs.apb_request_valid) {
                    data_state.apb.psel    <= 1;
                    data_state.apb.pwrite  <= (dmem_access_req.req_type == rv_mem_access_write);
                    data_state.apb.pwdata  <= dmem_access_req.write_data;
                    data_state.apb.paddr   <= dmem_access_req.address;
                }
            }
        }

        /*b APB request out */
        rv_apb_request = data_state.apb;

        /*b All done */
    }

    /*b RV APB targets */
    rv_apb_targets : {
        timer_apb_request = rv_apb_request;
        timer_apb_request.psel  = rv_apb_request.psel && (rv_apb_request.paddr[4;12]==0);
        timer_apb_request.paddr = rv_apb_request.paddr >> 2;

        apb_target_rv_timer tim( clk <- clk,
                                 reset_n <= reset_n,
                                 timer_control  <= timer_control,

                                 apb_request  <= timer_apb_request,
                                 apb_response => timer_apb_response,
                                 timer_value => timer_value );
        rv_apb_response = timer_apb_response;
    }

    /*b Instantiate debug
     */
    debug_instances: {
        tck_enable_fix = tck_enable;
        debug_tgt  = debug_tgt0;

        jtag_tap tap( jtag_tck <- jtag_tck_gated,
                      reset_n <= reset_n,
                      jtag <= jtag,
                      tdo => tdo,

                      ir => ir,
                      dr_action => dr_action,
                      dr_in => dr_in,
                      dr_tdi_mask <= dr_tdi_mask,
                      dr_out <= dr_out );

        riscv_jtag_apb_dm dm_apb( jtag_tck <- jtag_tck_gated,
                      reset_n <= reset_n,

                      ir <= ir,
                      dr_action <= dr_action,
                      dr_in <= dr_in,
                      dr_tdi_mask => dr_tdi_mask,
                      dr_out => dr_out,

                      apb_clock <- clk,
                      apb_request  => dm_apb_request,
                      apb_response <= dm_apb_response );

        riscv_i32_debug dm( clk <- clk,
                            reset_n <= reset_n,

                            apb_request  <= dm_apb_request,
                            apb_response => dm_apb_response,

                            debug_mst  => debug_mst,
                            debug_tgt <= debug_tgt 
            );
    }

    /*b Instantiate Reve-R pipeline
     */
    reve_r_pipeline: {
        riscv_i32_pipeline_control pc(clk <- clk,
                                      reset_n          <= reset_n,
                                      riscv_clk_enable <= riscv_clk_enable,
                                      csrs <= csrs,
                                      pipeline_state => pipeline_state,
                                      pipeline_response <= pipeline_response,
                                      pipeline_fetch_data <= pipeline_fetch_data,
                                      pipeline_control <= pipeline_control,
                                      riscv_config     <= riscv_config,
                                      trace            <= trace,
                                      debug_mst        <= debug_mst,
                                      debug_tgt       => debug_tgt0,
                                      rv_select <= 0 );

        riscv_i32_pipeline_control_fetch_req pc_fetch_req( pipeline_state <= pipeline_state,
                                                           pipeline_response <= pipeline_response,
                                                           pipeline_fetch_req => pipeline_fetch_req,
                                                           ifetch_req => rv_imem_access_req );

        riscv_i32_pipeline_control_fetch_data pc_fetch_data( pipeline_state <= pipeline_state,
                                                             ifetch_req  <= rv_imem_access_req,
                                                             ifetch_resp <= rv_imem_access_resp,
                                                             pipeline_fetch_req <= pipeline_fetch_req,
                                                             pipeline_fetch_data => pipeline_fetch_data );

        riscv_i32_pipeline_trap_interposer ti( pipeline_state         <= pipeline_state,
                                               pipeline_response      <= pipeline_response,
                                               dmem_access_resp       <= dmem_access_resp,
                                               pipeline_trap_request  => pipeline_trap_request,
                                               riscv_config           <= riscv_config
        );
        
        riscv_i32_pipeline_control_flow cf( pipeline_state <= pipeline_state,
                                            ifetch_req  <= rv_imem_access_req,
                                            pipeline_response <= pipeline_response,
                                            pipeline_trap_request  <= pipeline_trap_request,
                                            coproc_response <= coproc_response,
                                            pipeline_control => pipeline_control,
                                            dmem_access_resp <= dmem_access_resp,
                                            dmem_access_req => dmem_access_req,
                                            csr_access     => csr_access,
                                            pipeline_coproc_response => pipeline_coproc_response,
                                            coproc_controls  => coproc_controls,
                                            csr_controls     => csr_controls,
                                            trace            => trace,
                                            riscv_config <= riscv_config
        );
        
        riscv_i32c_pipeline3 dut( clk <- clk,
                                  reset_n <= reset_n,
                                  pipeline_control <= pipeline_control,
                                  pipeline_response => pipeline_response,
                                  pipeline_fetch_data <= pipeline_fetch_data,
                                  dmem_access_resp <= dmem_access_resp,
                                  coproc_response <= pipeline_coproc_response,
                                  csr_read_data    <= csr_data.read_data,
                                  riscv_config <= riscv_config);
        
    }

    /*b CSRs
     */
    csr_instance: {
        riscv_csrs_minimal csrs( clk <- clk,
                                 reset_n <= reset_n,
                                 riscv_clk_enable <= riscv_clk_enable,
                                 irqs <= irqs,
                                 csr_access     <= csr_access,
                                 csr_data       => csr_data,
                                 csr_controls   <= csr_controls,
                                 csrs => csrs
            );
    }
    
    /*b Coprocessors
     */
    coprocessors: {
        riscv_i32_muldiv m( clk <- clk,
                            reset_n <= reset_n,
                            coproc_controls <= coproc_controls,
                            coproc_response => coproc_response,
                            riscv_config <= riscv_config );

    }
    
    /*b Test harness
     */
    test_harness_inst: {
        se_test_harness th(clk <- jtag_tck, jtag=>jtag, tck_enable=>tck_enable, tdo<=tdo);
    }
    
    /*b Trace logic and modules
     */
    riscv_trace: {
        trace_control = {enable=1,
                         enable_control=1,
                         enable_pc=1, // priority over rfd?
                         enable_rfd=0,
                         enable_breakpoint=1,
                         valid = riscv_clk_enable};
        riscv_i32_trace trace(clk <- clk,
                              reset_n <= reset_n,
                              riscv_clk_enable <= riscv_clk_enable,
                              trace <= trace );
        riscv_i32_trace_pack trace_pack(clk <- clk,
                                        reset_n <= reset_n,
                                        trace_control <= trace_control,
                                        trace <= trace,
                                        packed_trace => packed_trace );
        riscv_i32_trace_compression trace_compression(packed_trace<=packed_trace,
                                                      compressed_trace => compressed_trace );
        riscv_i32_trace_decompression trace_decompression( compressed_nybbles <= compressed_trace.data,
                                                           decompressed_trace => decompressed_trace,
                                                           nybbles_consumed => nybbles_consumed );
    }

    /*b Checkers - for matching trace etc
     */
    checkers: {
        chk_riscv_ifetch checker_ifetch( clk <- clk,
                                         fetch_req <= rv_imem_access_req,
                                         fetch_resp <= rv_imem_access_resp
                                         //error_detected =>,
                                         //cycle => ,
            );
        chk_riscv_trace checker_trace( clk <- clk,
                                       trace <= trace
                                         //error_detected =>,
                                         //cycle => ,
            );
    }

    /*b All done
     */
}
