/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   riscv_csrs_minimal.cdl
 * @brief  Control/status registers for a minimal RISC-V implementation
 *
 * This file contains a module that implements the in-CPU CSRs
 * required by a RISC-V implementation.
 */

/*a Includes */
include "riscv_internal_types.h"

/*a Constants that can be overridden */
constant integer mimpid = 0;
constant integer misa = 0;
constant integer mvendorid = 0;
constant integer mhartid = 0;
constant integer mstatus = 0;

/*a Types */
/*t t_csr_write */
typedef struct {
    bit     enable     "Asserted if a CSR write is in progress";
    bit[32] data       "Write data, dependent on current CSR data potentially";
} t_csr_write;

/*a Module */
module riscv_csrs_minimal( clock clk                                   "RISC-V clock",
                           input bit reset_n                           "Active low reset",
                           input t_riscv_irqs          irqs            "Interrupts in to the CPU",
                           input t_riscv_csr_access    csr_access      "RISC-V CSR access, combinatorially decoded",
                           input t_riscv_word          csr_write_data  "Write data for the CSR access, later in the cycle than @csr_access possibly",
                           output t_riscv_csr_data     csr_data        "CSR respone (including read data), from the current @a csr_access",
                           input t_riscv_csr_controls  csr_controls    "Control signals to update the CSRs",
                           output t_riscv_csrs_minimal csrs            "CSR values"
    )
"""
This module implements a minimal set of RISC-V CSRs, as per v2.1 (May
2016) of the RISC-V instruction set manual user level ISA and v1.9.1
of the privilege architecture (Nov 2016), with the exception that
MTIME has been removed (as this seems to be the correct thing to do).

The privilege specifcation (v1.10) indicates:

* meip is read-only and is derived from the external irq in to this module

* mtip is read-only, cleared by writing to the memory-mapped timer comparator

* msip is read-write in a memory-mapped register somewhere

Hence the irqs structure must provide these three signals


Minimal CSRs as only machine mode and debug mode are supported.
In debug mode every register access is supported.
In machine mode then every register EXCEPT access to ??? is supported.

Given machine mode is the only mode supported:

* there are no SEI and UEI interrupt pins in to this module

* SEIP and UEIP are not supported

* STIP and UTIP are not supported

* SSIP and USIP are not supported

* mstatus.SIE and mstatus.UIE (and previous versions) are hardwired to 0

* mstatus.SPP and mstatus.UPP are hardwired to 0

The mip (machine interrupt pending register) therefore is:

{20b0, MEIP, 3b0, MTIP, 3b0, MSIP, 3b0}

The mie (machine interrupt enable register) is:

{20b0, MEIE, 3b0, MTIE, 3b0, MSIE, 3b0}


The instruction to the pipeline to request an interrupt (which is only
taken if an instruction is in uncommitted in the execution stage) must be generated using the
execution mode and the interrupt enable bits and the interrupt pending
bits.

Hence the 'take interrupt' is (mip & mie) != 0 && mstatus.MIE && (current mode >= machine mode) && (current mode != debug mode).

The required priority order is:

external interrupts, software interrupts, timer interrupts

If an instruction has been committed then it may trap, and the trap
will occur prior to an interrupt which happens after the commit
point. In this case there will be a trap, and the trapped instruction
will be fetched, and then an interrupt can be taken.

When an interrupt is taken the following occurs:

* MPP <= current execution mode (must be machine mode, as debug mode is not interruptible)

* mstatus.MPIE <= mstatus.MIE

Note that WFI should wait independent of mstatus.MIE for (mip & mie) != 0 (given machine mode only)
In debug mode WFI should be a NOP.

WFI may always be a NOP.

"""
{

    /*b State
     */
    default clock clk;
    default reset active_low reset_n;
    clocked t_riscv_csrs_minimal csrs={*=0};
    comb t_csr_write  csr_write;

    /*b CSR read/write
     */
    csr_read_write """
    CSR_ADDR_MSTATUS
    CSR_ADDR_MISA
    CSR_ADDR_MVENDORID
    CSR_ADDR_MARCHID
    CSR_ADDR_MIMPID
    CSR_ADDR_MHARTID
    """: {

        /*b Decode read data and 'illegal_access' for the CSR access */
        csr_data = {*=0};
        csr_data.illegal_access = 1;
        part_switch (csr_access.address) {
        case CSR_ADDR_CYCLE     : { csr_data.illegal_access=0; csr_data.read_data = csrs.cycles[32;0]; }
        case CSR_ADDR_CYCLEH    : { csr_data.illegal_access=0; csr_data.read_data = csrs.cycles[32;32]; }
        case CSR_ADDR_MCYCLE    : { csr_data.illegal_access=0; csr_data.read_data = csrs.cycles[32;0]; }
        case CSR_ADDR_MCYCLEH   : { csr_data.illegal_access=0; csr_data.read_data = csrs.cycles[32;32]; }
        case CSR_ADDR_INSTRET   : { csr_data.illegal_access=0; csr_data.read_data = csrs.instret[32;0]; }
        case CSR_ADDR_INSTRETH  : { csr_data.illegal_access=0; csr_data.read_data = csrs.instret[32;32]; }
        case CSR_ADDR_MINSTRET  : { csr_data.illegal_access=0; csr_data.read_data = csrs.instret[32;0]; }
        case CSR_ADDR_MINSTRETH : { csr_data.illegal_access=0; csr_data.read_data = csrs.instret[32;32]; }
        case CSR_ADDR_TIME      : { csr_data.illegal_access=0; csr_data.read_data = csrs.time[32;0]; }
        case CSR_ADDR_TIMEH     : { csr_data.illegal_access=0; csr_data.read_data = csrs.time[32;32]; }
        case CSR_ADDR_MIMPID    : { csr_data.illegal_access=0; csr_data.read_data = mimpid; }
        case CSR_ADDR_MHARTID   : { csr_data.illegal_access=0; csr_data.read_data = mhartid; }
        case CSR_ADDR_MISA      : { csr_data.illegal_access=0; csr_data.read_data = misa; }
        case CSR_ADDR_MVENDORID : { csr_data.illegal_access=0; csr_data.read_data = mvendorid; }
        case CSR_ADDR_MSTATUS   : { csr_data.illegal_access=0; csr_data.read_data = mstatus; }
        case CSR_ADDR_MSCRATCH  : { csr_data.illegal_access=0; csr_data.read_data = csrs.mscratch; }
        case CSR_ADDR_MEPC      : { csr_data.illegal_access=0; csr_data.read_data = csrs.mepc; }
        case CSR_ADDR_MCAUSE    : { csr_data.illegal_access=0; csr_data.read_data = csrs.mcause; }
        case CSR_ADDR_MTVAL     : { csr_data.illegal_access=0; csr_data.read_data = csrs.mtval; }
        case CSR_ADDR_MTVEC     : { csr_data.illegal_access=0; csr_data.read_data = csrs.mtvec; } // can be hardwired to any value, or read/write; tests require read-write
            // basic RISC-V tests require the following to not be illegal to write to
        case CSR_ADDR_MEDELEG   : { csr_data.illegal_access=0; csr_data.read_data = 0; } // must be 0 as only machine mode is supported
        case CSR_ADDR_MIDELEG   : { csr_data.illegal_access=0; csr_data.read_data = 0; } // must be 0 as only machine mode is supported
        case CSR_ADDR_MIE       : { csr_data.illegal_access=0; csr_data.read_data = 0; }
        }

        /*b Decode CSR writes */
        csr_write.enable = 0;
        csr_write.data = csr_write_data;
        part_switch (csr_access.access) {
        case riscv_csr_access_write: { csr_write.enable=1; }
        case riscv_csr_access_rw:    { csr_write.enable=1; }
        case riscv_csr_access_rs:    { csr_write.enable=1; csr_write.data |= csr_data.read_data; }
        case riscv_csr_access_rc:    { csr_write.enable=1; csr_write.data  = csr_data.read_data &~ csr_write_data; }
        }

        /*b All done */
    }

    /*b CSR state update */
    csr_state_update """
    """: {
        /*b Mirror time */
        csrs.time <= irqs.time;
            
        /*b Handle CSR cycle state */
        csrs.cycles[32;0] <= csrs.cycles[32;0] + 1;
        if (csrs.cycles[32;0]==-1) {csrs.cycles[32;32] <= csrs.cycles[32;32]+1;}

        if (csr_write.enable && (csr_access.address==CSR_ADDR_MCYCLE)) {
            csrs.cycles[32;0]    <= csr_write.data;
        }
        if (csr_write.enable && (csr_access.address==CSR_ADDR_MCYCLEH)) {
            csrs.cycles[32;32]    <= csr_write.data;
        }

        /*b Handle instruction retire counter state */
        if (csr_controls.retire) {
            csrs.instret[32;0] <= csrs.instret[32;0] + 1;
            if (csrs.instret[32;0]==-1) {csrs.instret[32;32] <= csrs.instret[32;32]+1;}
        }
        if (csr_write.enable && (csr_access.address==CSR_ADDR_MINSTRET)) {
            csrs.instret[32;0] <= csr_write.data;
        }
        if (csr_write.enable && (csr_access.address==CSR_ADDR_MINSTRETH)) {
            csrs.instret[32;32] <= csr_write.data;
        }

        /*b Handle MEPC state */
        if (csr_write.enable && (csr_access.address==CSR_ADDR_MEPC)) {
            csrs.mepc <= csr_write.data;
        }
        if (csr_controls.trap) {
            csrs.mepc <= csr_controls.trap_pc;
        }

        /*b Handle MTVEC state */
        if (csr_write.enable && (csr_access.address==CSR_ADDR_MTVEC)) {
            csrs.mtvec <= csr_write.data;
        }

        /*b Handle MTVAL state */
        if (csr_controls.trap) {
            csrs.mtval <= csr_controls.trap_value;
        }

        /*b Handle MCAUSE state */
        if (csr_write.enable && (csr_access.address==CSR_ADDR_MCAUSE)) {
            csrs.mcause <= csr_write.data;
        }
        if (csr_controls.trap) {
            full_switch (csr_controls.trap_cause) {
            case riscv_trap_cause_instruction_misaligned: { csrs.mcause <= bundle(24b0, riscv_mcause_instruction_misaligned); }
            case riscv_trap_cause_instruction_fault:      { csrs.mcause <= bundle(24b0, riscv_mcause_instruction_fault); }
            case riscv_trap_cause_illegal_instruction:    { csrs.mcause <= bundle(24b0, riscv_mcause_illegal_instruction); }
            case riscv_trap_cause_breakpoint:             { csrs.mcause <= bundle(24b0, riscv_mcause_breakpoint); }
            case riscv_trap_cause_load_misaligned:        { csrs.mcause <= bundle(24b0, riscv_mcause_load_misaligned); }
            case riscv_trap_cause_load_fault:             { csrs.mcause <= bundle(24b0, riscv_mcause_load_fault); }
            case riscv_trap_cause_store_misaligned:       { csrs.mcause <= bundle(24b0, riscv_mcause_store_misaligned); }
            case riscv_trap_cause_store_fault:            { csrs.mcause <= bundle(24b0, riscv_mcause_store_fault); }
            case riscv_trap_cause_uecall:                 { csrs.mcause <= bundle(24b0, riscv_mcause_uecall); }
            case riscv_trap_cause_secall:                 { csrs.mcause <= bundle(24b0, riscv_mcause_secall); }
            case riscv_trap_cause_hecall:                 { csrs.mcause <= bundle(24b0, riscv_mcause_hecall); }
            case riscv_trap_cause_mecall:                 { csrs.mcause <= bundle(24b0, riscv_mcause_mecall); }
            }
        }

        /*b Handle scratch state */
        if (csr_write.enable && (csr_access.address==CSR_ADDR_MSCRATCH)) {
            csrs.mscratch <= csr_write.data;
        }

        /*b All done */
    }

    /*b Logging */
    logging """
    """: {
        if (csr_write.enable) {
            if (csr_access.address == CSR_ADDR_DSCRATCH) {
                log("Scratch debug write",
                    "write_data", csr_write_data );
            }
        }
    }
}


