/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   riscv_minimal.cdl
 * @brief  Minimal RISC-V implementation ported to CDL
 *
 * CDL implementation of minimal RISC-V teaching implementation
 *
 * This is a two-stage pipeline implementation, with instruction fetch
 * of the next PC occuring simultaneously with the decode, register
 * read, ALU, data read/write request, data read memory access, and
 * register update.
 *
 * The instruction memory request, then, becomes valid dependent on
 * the decode of the registered instruction last fetched. For most
 * branches this requires only a small amount of logic, but for
 * jump-and-link-register instructions (which uses the full ALU
 * result) this may take a considerable amount of gates to determine
 * the correct branch target and hence next instruction fetch.  Hence
 * the instruction memory request is valid after a considerable delay
 * from the start of the cycle.
 *
 * The return value from the instruction memory request must be valid
 * before the end of the cycle.
 *
 * Any instruction memory implementation must start its access well
 * after the CPU clock edge, , as the request is valid after the CPU
 * clock edge; the resultant read data delay (from the clock edge)
 * then has to be factored in to determine when the next CPU clock
 * edge can occur. Hence it may be sensible to use a double speed
 * clock (e.g. 'fast_clk') to generate CPU clock edges (every other
 * fast_clk edge) and SRAM access clock edges (for a synchronous
 * memory) on the intervening fast_clk edges.
 *
 * The data memory request becomes valid, again, a fair time after the
 * CPU clock edge, as it requires instruction decode, register fetch,
 * and ALU operation to occur prior to the memory address being valid.
 *
 * The data memory response must be valid (for read data!) in the same
 * CPU cycle, as the returning data has to be rotated to the correct
 * byte lanes and prepared for the register file write.
 *
 * Hence a data memory implementation can be similar to that proposed
 * for the instruction memory - that is, accesses start on a memory
 * clock edge that is in the middle of a CPU clock edge, by using a
 * fast_clk.
 *
 */

/*a Includes
 */
include "cpu/riscv/riscv_internal_types.h"
include "cpu/riscv/riscv.h"
include "cpu/riscv/riscv_submodules.h"

/*a Constants
 */
constant integer INITIAL_PC=0x0;
constant integer i32c_force_disable=0;
constant integer coproc_force_disable=0;

/*a Types
 */
/*t t_decexecrfw_state */
typedef struct {
    t_riscv_i32_inst instruction   "Fetched instruction, ready for decode, register fetch, execute and writeback";
    bit valid                      "Asserted if @instr_data is a valid fetched instruction, whether misaligned or not";
    bit[32] pc                     "PC of the fetched instruction";
} t_decexecrfw_state;

/*t t_decexecrfw_combs
 *
 * Combinatorials of the decexecrfw_state
 */
typedef struct {
    t_riscv_i32_decode idecode;

    t_riscv_word   rs1;
    t_riscv_word   rs2;

    bit exec_committed;
    t_riscv_csr_access csr_access;
    t_riscv_word rfw_write_data;
    t_riscv_i32_dmem_exec dmem_exec;
    t_riscv_i32_control_data control_data;
} t_decexecrfw_combs;

/*a Module
 */
module riscv_i32c_pipeline( clock clk,
                            input bit reset_n,
                            input t_riscv_irqs       irqs               "Interrupts in to the CPU",
                            output t_riscv_mem_access_req      dmem_access_req,
                            input  t_riscv_mem_access_resp     dmem_access_resp,
                            input t_riscv_pipeline_control     pipeline_control,
                            output t_riscv_pipeline_response   pipeline_response,
                            input t_riscv_pipeline_fetch_data  pipeline_fetch_data,
                            output t_riscv_i32_coproc_controls coproc_controls,
                            input t_riscv_i32_coproc_response  coproc_response,
                            input  t_riscv_config              riscv_config,
                            output t_riscv_csrs_minimal        csrs,
                            output t_riscv_i32_trace           trace
)
"""
This is just the processor pipeline, using a single stage for execution.

The instruction fetch request for the next cycle is put out just after
the ALU stage logic, which may be a long time into the cycle; the
fetch data response presents the instruction fetched at the end of the
cycle, where it is registered for execution.

The pipeline is then a single stage that takes the fetched
instruction, decodes, fetches register values, and executes the ALU
stage; determining in half a cycle the next instruction fetch, and in
the whole cycle the data memory request, which is valid just before
the end

A coprocessor is supported; this may be configured to be disabled, in
which case the outputs are driven low and the inputs are coprocessor
response is ignored.

A coprocessor can implement, for example, the multiply for i32m (using
riscv_i32_muldiv).  Note that since there is not a separate decode
stage the multiply cannot support fused operations

"""
{

    /*b State and comb
     */
    default clock clk;
    default reset active_low reset_n;

    clocked t_riscv_word[32] registers={*=0} "Register 0 is tied to 0 - so it is written on every cycle to zero...";

    net     t_riscv_i32_decode     decexecrfw_idecode_i32;
    net     t_riscv_i32_decode     decexecrfw_idecode_i32c;
    clocked t_decexecrfw_state     decexecrfw_state={*=0, pc=INITIAL_PC};
    comb    t_decexecrfw_combs     decexecrfw_combs;
    net     t_riscv_i32_dmem_request decexecrfw_dmem_request "Data memory request data";
    net     t_riscv_word           decexecrfw_dmem_read_data;
    net     t_riscv_i32_control_flow decexecrfw_control_flow;
    net     t_riscv_i32_alu_result decexecrfw_alu_result;

    comb t_riscv_csr_controls csr_controls;
    net t_riscv_csr_data csr_data;
    net t_riscv_csrs_minimal csrs;

    /*b Decode, RFR, execute and RFW stage - single stage execution
     */
    decode_rfr_execute_stage """
    The decode/RFR/execute stage performs all of the hard workin the
    implementation.

    It first incorporates a program counter (PC) and an instruction
    register (IR). The instruction in the IR corresponds to that
    PC. Initially (at reset) the IR will not be valid, as an
    instruction must first be fetched, so there is a corresponding
    valid bit too.

    The IR is decoded as both a RV32C (16-bit) and RV32 (32-bit) in
    parallel; the bottom two bits of the instruction register indicate
    which is valid for the IR.

    """: {
        /*b Instruction register - note all PC value are legal (bit 0 is cleared automatically though) */
        decexecrfw_state.valid <= 0;
        if (pipeline_fetch_data.valid) {
            decexecrfw_state.instruction <= {
                data = pipeline_fetch_data.data,
                mode = pipeline_control.mode };
            decexecrfw_state.valid <= 1;
            decexecrfw_state.pc <= pipeline_fetch_data.pc;
        }

        /*b Decode instruction */
        riscv_i32_decode decode_i32( instruction <= decexecrfw_state.instruction,
                                     idecode      => decexecrfw_idecode_i32,
                                     riscv_config <= riscv_config );

        riscv_i32c_decode decode_i32c( instruction <= decexecrfw_state.instruction,
                                       idecode      => decexecrfw_idecode_i32c,
                                       riscv_config <= riscv_config );

        /*b Select decode (from either i32 or i32c or possible debug) */
        decexecrfw_combs.idecode = decexecrfw_idecode_i32;
        if ((!i32c_force_disable) && riscv_config.i32c) {
            if (decexecrfw_state.instruction.data[2;0]!=2b11) {
                decexecrfw_combs.idecode = decexecrfw_idecode_i32c;
            }
        }

        /*b Determine whether to commit to execute */
        decexecrfw_combs.exec_committed = decexecrfw_state.valid;
        if (decexecrfw_combs.idecode.illegal || decexecrfw_combs.idecode.illegal_pc) {
            decexecrfw_combs.exec_committed = 0;
        }
        // block interrupt_req if in second+ cycle of multicycle exec operation
        if (pipeline_control.interrupt_req) {
            decexecrfw_combs.exec_committed = 0;
        }

        /*b Register read - post decode, prior to ALU and CSRs */
        decexecrfw_combs.rs1 = registers[decexecrfw_combs.idecode.rs1]; // note that register 0 is ALWAYS 0 anyway
        decexecrfw_combs.rs2 = registers[decexecrfw_combs.idecode.rs2]; // note that register 0 is ALWAYS 0 anyway

        /*b Execute ALU stage - post register read, parallel with CSRs */
        riscv_i32_alu alu( idecode <= decexecrfw_combs.idecode,
                           pc  <= decexecrfw_state.pc,
                           rs1 <= decexecrfw_combs.rs1,
                           rs2 <= decexecrfw_combs.rs2,
                           alu_result => decexecrfw_alu_result );
    
        /*b Minimal CSRs - post register read, parallel with ALU */
        decexecrfw_combs.csr_access                  = decexecrfw_combs.idecode.csr_access;
        decexecrfw_combs.csr_access.access_cancelled = !decexecrfw_combs.exec_committed;
        decexecrfw_combs.csr_access.write_data       = decexecrfw_combs.idecode.immediate_valid ? bundle(27b0, decexecrfw_combs.idecode.rs1) : decexecrfw_combs.rs1;
        riscv_csrs_minimal csrs( clk <- clk,
                                 reset_n <= reset_n,
                                 irqs <= irqs,
                                 csr_access     <= decexecrfw_combs.csr_access,
                                 csr_data       => csr_data,
                                 csr_controls   <= csr_controls,
                                 csrs => csrs);

        /*b Memory access handling - post ALU - must be valid before middle of cycle */
        decexecrfw_combs.dmem_exec = { idecode = decexecrfw_combs.idecode,
                                       arith_result   = decexecrfw_alu_result.arith_result, // address of access
                                       rs2            = decexecrfw_combs.rs2,    // data for access (before rotation)
                                       exec_committed = decexecrfw_combs.exec_committed,
                                       first_cycle = 1
        };
        riscv_i32_dmem_request dmem_req( dmem_exec    <= decexecrfw_combs.dmem_exec,
                                         dmem_request => decexecrfw_dmem_request );
        dmem_access_req = decexecrfw_dmem_request.access;
        // should use illegal dmem access for trap
        // should use 'needs second cycle'

        /*b Control flow - post ALU for next PC & branch condition met, rest from decode */
        decexecrfw_combs.control_data = { instruction_data = decexecrfw_state.instruction.data,
                                          pc = decexecrfw_state.pc,
                                          alu_result = decexecrfw_alu_result,
                                          interrupt_ack = 1,
                                          exec_committed = decexecrfw_combs.exec_committed,
                                          idecode = decexecrfw_combs.idecode,
                                          first_cycle = 1
        };
        riscv_i32_control_flow control_flow( pipeline_control <= pipeline_control,
                                             control_data <= decexecrfw_combs.control_data,
                                             control_flow => decexecrfw_control_flow );

        /*b Pipeline response from decode */
        // possible add in valid and illegal (if valid && illegal then pipeline will flush)
        pipeline_response.decode.valid         = decexecrfw_state.valid;
        pipeline_response.decode.pc            = decexecrfw_state.pc;
        pipeline_response.decode.is_compressed = decexecrfw_combs.idecode.is_compressed;
        pipeline_response.decode.action        = rv_pipe_dpc_sequential;
        pipeline_response.decode.branch_target = decexecrfw_alu_result.branch_target; // used only if predict_branch - i.e. never in this pipeline

        /*b Pipeline response from exec */
        pipeline_response.exec.valid = decexecrfw_state.valid;
        pipeline_response.exec.interrupt_ack = pipeline_control.interrupt_req;
        pipeline_response.exec.trap = {*=0};
        pipeline_response.exec.is_compressed = decexecrfw_combs.idecode.is_compressed;
        pipeline_response.exec.pc            = decexecrfw_state.pc;
        pipeline_response.exec.action        = rv_pipe_epc_predicted; // Normal action is Exec follows whatever was decoded (if there was anything)
        pipeline_response.exec.flush_target = decexecrfw_alu_result.branch_target;

        if (decexecrfw_control_flow.branch_taken) {
            pipeline_response.exec.action = rv_pipe_epc_flush;
        }
        pipeline_response.exec.trap = decexecrfw_control_flow.trap;

        /*b CSR controls - post trap detection */
        csr_controls = {*=0};
        csr_controls.retire       = decexecrfw_combs.exec_committed;
        csr_controls.trap         = decexecrfw_control_flow.trap;
        csr_controls.trap.to_mode = rv_mode_machine;

        /*b Memory read handling - post memory request and memory read - so way late in the second half of the cycle */
        riscv_i32_dmem_read_data dmem_data( dmem_request <= decexecrfw_dmem_request,
                                            last_data <= 0, // only for unaligned reads
                                            dmem_access_resp <= dmem_access_resp,
                                            dmem_read_data => decexecrfw_dmem_read_data);

        /*b Register write - post memory read
         */
        decexecrfw_combs.rfw_write_data = decexecrfw_alu_result.result | coproc_response.result;
        if (coproc_force_disable || riscv_config.coproc_disable) {
            decexecrfw_combs.rfw_write_data = decexecrfw_alu_result.result;
        }
        if (dmem_access_req.read_enable) {
            decexecrfw_combs.rfw_write_data =  decexecrfw_dmem_read_data;
        }
        if (decexecrfw_combs.idecode.csr_access.access != riscv_csr_access_none) {
            decexecrfw_combs.rfw_write_data = csr_data.read_data;
        }
        if (decexecrfw_combs.exec_committed && decexecrfw_combs.idecode.rd_written) {
            registers[decexecrfw_combs.idecode.rd] <= decexecrfw_combs.rfw_write_data;
        }
        registers[0] <= 0; // register 0 is always zero...
    }

    /*b Coprocessor interface */
    coprocessor_interface """
    Drive the coprocessor controls unless disabled; mirror the pipeline combs
    """: {
        coproc_controls = {*=0};
        coproc_controls.dec_idecode_valid  = decexecrfw_state.valid && !pipeline_control.interrupt_req;
        coproc_controls.dec_idecode        = decexecrfw_combs.idecode;
        coproc_controls.dec_to_alu_blocked = coproc_response.cannot_complete; // If ALU can complete...
        coproc_controls.alu_rs1 = decexecrfw_combs.rs1;
        coproc_controls.alu_rs2 = decexecrfw_combs.rs2;
        coproc_controls.alu_flush_pipeline = 0; // No pipeline to flush
        coproc_controls.alu_cannot_start = coproc_response.cannot_start;       // ALU can always start itself; coprocessor can block it
        coproc_controls.alu_cannot_complete = coproc_response.cannot_complete; // ALU can always complete (no unaligned transactions yet); coprocessor can block it
        if (coproc_force_disable || riscv_config.coproc_disable) {
            coproc_controls = {*=0};
        }
    }

    /*b Logging */
    logging """
    """: {
        trace = {*=0};
        trace.instr_valid    = decexecrfw_combs.exec_committed;
        trace.instr_pc       = pipeline_response.exec.pc;
        trace.instruction    = decexecrfw_state.instruction;
        trace.rfw_retire     = csr_controls.retire;
        trace.rfw_data_valid = decexecrfw_combs.idecode.rd_written && decexecrfw_combs.exec_committed;
        trace.rfw_rd         = decexecrfw_combs.idecode.rd;
        trace.rfw_data       = decexecrfw_combs.rfw_write_data;
        trace.branch_taken   = decexecrfw_control_flow.branch_taken;
        trace.trap           = decexecrfw_control_flow.trap.valid;
        trace.branch_target  = pipeline_response.exec.flush_target;
    }

    /*b All done */
}

