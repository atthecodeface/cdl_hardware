/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   riscv_minimal.cdl
 * @brief  Minimal RISC-V implementation ported to CDL
 *
 * CDL implementation of minimal RISC-V teaching implementation
 *
 * This is a two-stage pipeline implementation, with instruction fetch
 * of the next PC occuring simultaneously with the decode, register
 * read, ALU, data read/write request, data read memory access, and
 * register update.
 *
 * The instruction memory request, then, becomes valid dependent on
 * the decode of the registered instruction last fetched. For most
 * branches this requires only a small amount of logic, but for
 * jump-and-link-register instructions (which uses the full ALU
 * result) this may take a considerable amount of gates to determine
 * the correct branch target and hence next instruction fetch.  Hence
 * the instruction memory request is valid after a considerable delay
 * from the start of the cycle.
 *
 * The return value from the instruction memory request must be valid
 * before the end of the cycle.
 *
 * Any instruction memory implementation must start its access well
 * after the CPU clock edge, , as the request is valid after the CPU
 * clock edge; the resultant read data delay (from the clock edge)
 * then has to be factored in to determine when the next CPU clock
 * edge can occur. Hence it may be sensible to use a double speed
 * clock (e.g. 'fast_clk') to generate CPU clock edges (every other
 * fast_clk edge) and SRAM access clock edges (for a synchronous
 * memory) on the intervening fast_clk edges.
 *
 * The data memory request becomes valid, again, a fair time after the
 * CPU clock edge, as it requires instruction decode, register fetch,
 * and ALU operation to occur prior to the memory address being valid.
 *
 * The data memory response must be valid (for read data!) in the same
 * CPU cycle, as the returning data has to be rotated to the correct
 * byte lanes and prepared for the register file write.
 *
 * Hence a data memory implementation can be similar to that proposed
 * for the instruction memory - that is, accesses start on a memory
 * clock edge that is in the middle of a CPU clock edge, by using a
 * fast_clk.
 *
 */

/*a Includes
 */
include "cpu/riscv/riscv.h"
include "cpu/riscv/riscv_modules.h"

/*a Module
 */
module riscv_i32_minimal_apb( clock clk,
                              input bit reset_n,
                              input  t_riscv_mem_access_req  data_access_req,
                              output t_riscv_mem_access_resp data_access_resp,
                              output t_apb_request apb_request,
                              input  t_apb_response apb_response
)
"""
"""
{

    /*b State and comb
     */
    default clock clk;
    default reset active_low reset_n;
    clocked t_apb_request apb_request={*=0};

    apb_logic "": {
        data_access_resp = {*=0};
        data_access_resp.ack = 1;
        data_access_resp.ack_if_seq = 1;
        data_access_resp.abort_req = 0;
        data_access_resp.access_complete = 1;
        if (apb_request.penable) {
            data_access_resp.read_data = apb_response.prdata;
        }

        if (apb_request.psel) {
            data_access_resp.ack = 0;
            data_access_resp.ack_if_seq = 0;
            data_access_resp.access_complete = 0;
            apb_request.penable <= 1;
            if (apb_request.penable && apb_response.pready) {
                apb_request.psel <= 0;
                apb_request.penable <= 0;
                data_access_resp.access_complete = 1;
            }
        } else {
            if (data_access_req.valid) {
                apb_request.psel <= 1;
                apb_request.penable <= 0;
                apb_request.paddr <= data_access_req.address;
                apb_request.pwrite <= (data_access_req.req_type == rv_mem_access_write);
                apb_request.pwdata <= data_access_req.write_data;
            }
        }
    }
}
