/** @copyright (C) 2020,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   teletext_dprintf_mux.cdl
 * @brief  A valid/ack multiplexer to dprintf requests
 *
 * Use of the generic utility valid/ack multiplexer
 *
 * Needs to be built in CDL with the options:
 *
 *  rmt:gt_generic_valid_req=t_dprintf_req_4
 *
 *  rmn:generic_valid_fifo=dprintf_4_fifo
 *
 *  dc:fifo_depth=3
 *
 * The FIFO depth in the constant can be 1 less than the required size as the FIFO as an output register
 */
/*a Includes */
include "types/dprintf.h"

/*a Module */
include "generic_valid_ack_sram_fifo.cdl"
