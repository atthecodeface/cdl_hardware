/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   tb_kasumi_cipher.cdl
 * @brief  Testbench for Kasumi cipher modules
 *
 */

/*a Includes
 */
include "crypt/kasumi_types.h"
include "crypt/kasumi_modules.h"

/*a External modules */
extern module se_test_harness( clock clk, output t_kasumi_input kasumi_input, input bit kasumi_input_ack, input t_kasumi_output kasumi_output, output bit kasumi_output_ack )
{
    timing from rising clock clk kasumi_input, kasumi_output_ack;
    timing to   rising clock clk kasumi_output, kasumi_input_ack;
}

/*a Module
 */
module tb_kasumi_cipher( clock clk,
                         input bit reset_n
)
{

    /*b Nets
     */
    net t_kasumi_input    kasumi_input;
    net bit              kasumi_input_ack;
    net t_kasumi_output  kasumi_output;
    net bit               kasumi_output_ack;

    /*b Instantiate RISC-V
     */
    riscv_instance: {
        se_test_harness th( clk <- clk,
                            kasumi_input => kasumi_input,
                            kasumi_output_ack => kasumi_output_ack,

                            kasumi_input_ack <= kasumi_input_ack,
                            kasumi_output    <= kasumi_output );
        
        kasumi_cipher dut(   clk <- clk,
                             reset_n <= reset_n,
                             kasumi_input_ack => kasumi_input_ack,
                             kasumi_output    => kasumi_output,
                             kasumi_input <= kasumi_input,
                             kasumi_output_ack <= kasumi_output_ack );

    }
}
