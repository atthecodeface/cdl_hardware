/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   dprintf.cdl
 * @brief  Debug text formatter
 *
 * CDL implementation of a module that takes an input debug requests
 * and converts them in to a stream of bytes. The debug request is
 * similar to a 'printf' string, in that it allows formatted data.
 *
 */
/*a Includes */
include "srams.h"
include "types/dprintf.h"

/*a Module
 */
module dprintf_4_dp_sram_512(
    clock write_clk,
    clock read_clk,
    input bit write_enable,
    input bit[9] write_address,
    input t_dprintf_req_4 write_data,
    input bit read_enable,
    input bit[9] read_address,
    output t_dprintf_req_4 read_data
    )
"""
Map dprintf_4 to dual-port SRAMs.
"""
{
    comb bit[64][4] sr_write_data;
    net bit[32]     sr_read_address;
    net bit[64][4]  sr_read_data;
    srams: {
        se_sram_mrw_2_512x32 sr_ctl( sram_clock_0 <- write_clk,
                                     select_0 <= write_enable,
                                     address_0 <= write_address,
                                     read_not_write_0 <= 0,
                                     // data_out_0,
                                     sram_clock_1 <- read_clk,
                                     select_1 <= read_enable,
                                     address_1 <= read_address,
                                     read_not_write_1 <= 1,
                                     write_data_1 <= 0,

                                     write_data_0 <= bundle(16b0, write_data.address),
                                     data_out_1 => sr_read_address
            );
        for (i; 4) {
            se_sram_mrw_2_512x64 sr_data[i]( sram_clock_0 <- write_clk,
                                             select_0 <= write_enable,
                                             address_0 <= write_address,
                                             read_not_write_0 <= 0,
                                             // data_out_0,
                                             sram_clock_1 <- read_clk,
                                             select_1 <= read_enable,
                                             address_1 <= read_address,
                                             read_not_write_1 <= 1,
                                             write_data_1 <= 0,

                                             write_data_0 <= sr_write_data[i],
                                             data_out_1 => sr_read_data[i]
                );
        }
        sr_write_data[0] = write_data.data_0;
        sr_write_data[1] = write_data.data_1;
        sr_write_data[2] = write_data.data_2;
        sr_write_data[3] = write_data.data_3;
        read_data.valid = 0;
        read_data.address = sr_read_address[16;0];
        read_data.data_0 = sr_read_data[0];
        read_data.data_1 = sr_read_data[1];
        read_data.data_2 = sr_read_data[2];
        read_data.data_3 = sr_read_data[3];
    }
}
