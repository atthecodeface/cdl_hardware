/** @copyright (C) 2019,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   apb_target_uart_minimal.cdl
 * @brief  A minimal UART with single tx/rx holding bytes
 *
 * CDL implementation of a very simple APB UART
 */
/*a Includes */
include "types/apb.h"
include "types/uart.h"
include "types/clock_divider.h"
include "input/uart_modules.h"
include "utils/clock_divider_modules.h"

/*a Constants
*/

/*a Types
*/
/*t t_apb_access - Read or write action due to APB request */
typedef enum[4] {
    apb_access_none,
    apb_access_write_config,
    apb_access_read_config,
    apb_access_write_brg,
    apb_access_read_brg,
    apb_access_write_holding,
    apb_access_read_holding,
    apb_access_read_status
} t_apb_access;

/*t t_apb_state - clocked state for APB side */
typedef struct {
    t_apb_access access;
} t_apb_state;

/*t t_apb_address */
typedef enum[3] {
    apb_address_status  = 0,
    apb_address_brg     = 1,
    apb_address_config  = 2,
    apb_address_holding = 3
} t_apb_address;

/*a Module
*/
/*m apb_target_uart_minimal */
module apb_target_uart_minimal( clock clk,
                                input bit reset_n,

                                input  t_apb_request  apb_request  "APB request",
                                output t_apb_response apb_response "APB response",

                                input    t_uart_rx_data uart_rx,
                                output   t_uart_tx_data uart_tx,
                                output   t_uart_status  status
    )
"""
This is an APB target that uses a minimal UART
"""
{
    /*b Default clock/reset */
    default clock clk;
    default reset active_low reset_n;

    /*b APB interface state  */
    clocked t_apb_state    apb_state   = {*=0}  "Decode of APB";

    /*b UART signals */
    comb t_uart_control uart_control;
    net t_uart_output   uart_output;
    net t_uart_tx_data  uart_tx;
    
    /*b Outputs */
    drive_outputs : {
        status = uart_output.status;
    }

    /*b APB interface */
    apb_interface : {

        /*b APB interface decode */
        part_switch (apb_request.paddr[3;0]) {
        case apb_address_status: {
            apb_state.access  <= apb_request.pwrite ? apb_access_none : apb_access_read_status;
        }
        case apb_address_config: {
            apb_state.access  <= apb_request.pwrite ? apb_access_write_config : apb_access_read_config;
        }
        case apb_address_brg: {
            apb_state.access  <= apb_request.pwrite ? apb_access_write_brg : apb_access_read_brg;
        }
        case apb_address_holding: {
            apb_state.access  <= apb_request.pwrite ? apb_access_write_holding : apb_access_read_holding;
        }
        }
        if (!apb_request.psel || apb_request.penable) {
            apb_state.access <= apb_access_none;
        }

        /*b APB interface response - use apb_state.access */
        apb_response = {*=0, pready=1};
        part_switch (apb_state.access) {
        case apb_access_read_status: {
            apb_response.prdata[8]  = !uart_output.tx_ack;
            apb_response.prdata[16] = uart_output.rx_valid;
            apb_response.prdata[17] = uart_output.status.rx_half_full;
            apb_response.prdata[18] = uart_output.status.rx_overflow;
            apb_response.prdata[19] = uart_output.status.rx_framing_error;
            apb_response.prdata[20] = uart_output.status.rx_parity_error;
        }
        case apb_access_read_config: {
            apb_response.prdata = uart_output.config_data;
        }
        case apb_access_read_brg: {
            apb_response.prdata = uart_output.brg_config_data;
        }
        case apb_access_read_holding: {
            apb_response.prdata[8;0] = uart_output.rx_data;
            apb_response.prdata[28]  = uart_output.status.rx_overflow;
            apb_response.prdata[29]  = uart_output.status.rx_framing_error;
            apb_response.prdata[30]  = uart_output.status.rx_parity_error;
            apb_response.prdata[31]  = !uart_output.rx_valid;
        }
        }

        /*b All done */
    }
        
    /*b UART instance */
    uart_instance """
    """ : {
        uart_control.clear_errors = (apb_state.access==apb_access_read_status);
        uart_control.rx_ack       = (apb_state.access==apb_access_read_holding);
        uart_control.tx_valid     = (apb_state.access==apb_access_write_holding);
        uart_control.tx_data      = apb_request.pwdata[8;0];
        uart_control.write_config = (apb_state.access==apb_access_write_config);
        uart_control.write_brg    = (apb_state.access==apb_access_write_brg);
        uart_control.write_data   = apb_request.pwdata;

        uart_minimal uart(clk <- clk,
                          reset_n <= reset_n,
                          uart_control <= uart_control,
                          uart_output  => uart_output,
                          uart_rx <= uart_rx,
                          uart_tx => uart_tx );

        /*b All done */
    }

    /*b All done */
}
