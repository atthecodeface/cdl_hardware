/** @copyright (C) 2018,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   tb_riscv_jtag_debug.cdl
 * @brief  Testbench for RISC-V debug over JTAG
 *
 */

/*a Includes
 */
include "types/jtag.h"
include "types/apb.h"
include "cpu/riscv/riscv.h"
include "cpu/riscv/riscv_pipeline_types.h"
include "cpu/riscv/riscv_pipeline.h"
include "cpu/riscv/riscv_modules.h"

/*a External modules */
extern module se_test_harness( clock clk, output t_jtag jtag, output bit tck_enable, input bit tdo )
{
    timing from rising clock clk jtag, tck_enable;
    timing to rising clock clk tdo;
}

typedef struct {
    bit running;
    bit halting;
    bit resuming;
    bit resumed;
    bit attention;
    bit[8] counter;
} t_test_state;

/*a Module
 */
module tb_riscv_jtag_debug( clock jtag_tck,
                          clock apb_clock,
                          input bit reset_n
)
{

    /*b Nets
     */
    net t_jtag jtag;
    net bit tdo;
    net bit[5]ir;
    net t_jtag_action dr_action;
    net bit[50]dr_in;
    net bit[50]dr_tdi_mask;
    net bit[50]dr_out;
    net bit tck_enable;
    comb bit tck_enable_fix;
    gated_clock clock jtag_tck active_high tck_enable_fix jtag_tck_gated;

    net   t_apb_request  apb_request  "APB request";
    net   t_apb_response apb_response "APB response";
    net   t_riscv_debug_mst debug_mst;
    comb  t_riscv_debug_tgt debug_tgt;
    net   t_riscv_debug_tgt debug_tgt0;
    net   t_riscv_debug_tgt debug_tgt1;

    /*b Instantiate APB timer
     */
    net t_riscv_pipeline_state     pipeline_state0;
    net t_riscv_pipeline_state     pipeline_state1;
    comb t_riscv_pipeline_response   pipeline_response;
    comb t_riscv_pipeline_fetch_data  pipeline_fetch_data;
    comb t_riscv_i32_trace trace;
    comb t_riscv_csrs_minimal csrs;
    comb t_riscv_config riscv_config;
    dut_instance: {
        tck_enable_fix = tck_enable;
        riscv_config = {*=0};
        riscv_config.debug_enable = 1;
        pipeline_response = {*=0};
        pipeline_fetch_data = {*=0};
        trace = {*=0};
        csrs = {*=0};
        debug_tgt  = debug_tgt0;
        debug_tgt |= debug_tgt1;
        se_test_harness th(clk <- jtag_tck, jtag=>jtag, tck_enable=>tck_enable, tdo<=tdo);

        jtag_tap tap( jtag_tck <- jtag_tck_gated,
                      reset_n <= reset_n,
                      jtag <= jtag,
                      tdo => tdo,

                      ir => ir,
                      dr_action => dr_action,
                      dr_in => dr_in,
                      dr_tdi_mask <= dr_tdi_mask,
                      dr_out <= dr_out );

        riscv_jtag_apb_dm dm_apb( jtag_tck <- jtag_tck_gated,
                      reset_n <= reset_n,

                      ir <= ir,
                      dr_action <= dr_action,
                      dr_in <= dr_in,
                      dr_tdi_mask => dr_tdi_mask,
                      dr_out => dr_out,

                      apb_clock <- apb_clock,
                      apb_request => apb_request,
                      apb_response <= apb_response );

        riscv_i32_debug dm( clk <- apb_clock,
                            reset_n <= reset_n,

                            apb_request <= apb_request,
                            apb_response => apb_response,

                            debug_mst  => debug_mst,
                            debug_tgt <= debug_tgt 
            );
        riscv_i32_pipeline_control pc0(clk <- apb_clock,
                                                 reset_n <= reset_n,
                                       riscv_clk_enable <= 1,
                                                 csrs <= csrs,
                                                 pipeline_state => pipeline_state0,
                                                 pipeline_response <= pipeline_response,
                                                 pipeline_fetch_data <= pipeline_fetch_data,
                                                 riscv_config     <= riscv_config,
                                                 trace            <= trace,
                                                 debug_mst        <= debug_mst,
                                                 debug_tgt       => debug_tgt0,
                                                 rv_select <= 0 );
        riscv_i32_pipeline_control pc1(clk <- apb_clock,
                                                 reset_n <= reset_n,
                                       riscv_clk_enable <= 1,
                                                 csrs                <= csrs,
                                                 pipeline_state    => pipeline_state1,
                                                 pipeline_response   <= pipeline_response,
                                                 pipeline_fetch_data <= pipeline_fetch_data,
                                                 riscv_config        <= riscv_config,
                                                 trace               <= trace,
                                                 debug_mst           <= debug_mst,
                                                 debug_tgt           => debug_tgt1,
                                                 rv_select <= 1 );
    }
}
