/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   riscv_i32_alu.cdl
 * @brief  ALU for i32 RISC-V implementation
 *
 * CDL implementation of RISC-V i32 ALU based on the RISC-V
 * specification v2.1.
 *
 */

/*a Includes
 */
include "cpu/riscv/riscv_config.h"
include "cpu/riscv/riscv_internal_types.h"
include "cpu/riscv/riscv.h"

/*a Types
 */
/*t t_mask_type */
typedef enum[2] {
    mask_type_none    = 2b00,
    mask_type_normal  = 2b01,
    mask_type_invert  = 2b11,
    mask_type_rs2     = 2b10,
} t_mask_type;

/*t t_bbmask_type */
typedef enum[2] {
    bb_mask_type_all   = 2b00,
    bb_mask_type_bit   = 2b01,
    bb_mask_type_byte     = 2b11,
} t_bb_mask_type;

/*t t_shift_combs */
typedef struct {
    t_mask_type and_mask_type;
    t_mask_type or_mask_type;
    t_bb_mask_type bb_mask_type;
    bit[5]  shift_control;
    bit[5]  shift_amount;
    bit[32] rotate_in           "Data to rotate";
    bit[32] rotate_by_16        "Rotated optionally by 16";
    bit[32] rotate_byte_reverse "Optional byte reverse of rotate_by_16";
    bit[32] rotate_bit_reverse  "Optional bit reverse of rotate_byte_reverse";
    bit[48] rotate_out          "Bottom 32 bits only are used; this is rotate_by_16 duplicated >> (0 to 15)";
    bit[64] mask_in;
    bit[64] mask_out;
    bit[32] shift_and_mask;
    bit[32] shift_or_mask;
    bit[32] shift_result "Only bottom 32 bits are used";
} t_shift_combs;

/*t t_alu_combs */
typedef struct {
    t_riscv_word  imm_or_rs2;
    t_riscv_word  imm_or_rs1;
    bit[32] arith_in_0;
    bit[32] arith_in_1;
    bit     arith_carry_in;
    bit     carry_in_to_31;
    bit[32] arith_result_32;
    bit[33] arith_result;
    bit     arith_eq;
    bit     arith_unsigned_ge;
    bit     arith_signed_ge;
    t_riscv_word  pc_plus_4;
    t_riscv_word  pc_plus_2;
    t_riscv_word  pc_plus_inst;
    t_riscv_word  pc_plus_imm;
} t_alu_combs;

/*a Module
 */
module riscv_i32_alu( input t_riscv_i32_decode      idecode,
                      input t_riscv_word            pc,
                      input t_riscv_word            rs1,
                      input t_riscv_word            rs2,
                      output t_riscv_i32_alu_result alu_result
)
"""

"""
{

    /*b Signals - just the combs */
    comb t_shift_combs shift_combs    "Combinatorials used in the shifter";
    comb t_alu_combs   alu_combs      "Combinatorials used in the module, not exported as the decode";

    /*b Shifter operation */
    shifter_operation """
    The shifter can be built as a 64-bit shift-right-by-N, with masks to combine the two halves


    A rotate right by 
    """ : {
        shift_combs.and_mask_type = mask_type_none; // values for rotate (why not?)
        shift_combs.or_mask_type  = mask_type_none;
        shift_combs.bb_mask_type  = bb_mask_type_all;

        /*b Decode shift op
          Mask is ffff0000 >> amount
          shift left logical of zeros is (rotate and mask)
          shift left logical of ones is (rotate and mask) OR (~mask)
          shift right logical of zeros is (rotate and ~mask)
          shift right logical of ones is (rotate and ~mask) OR (mask)
          shift right arithmetic is (rotate and ~mask) OR ([31]?mask:0)
          rotate right/left is rotate
          reverse is reverse output

constant integer rv_cfg_i32_bitmap_enhanced_shift_enable=0;
constant integer rv_cfg_i32_bitmap_others_enable=0;

         */
        part_switch (idecode.shift_op) {
        case riscv_shift_op_left_logical_zeros:   {
            shift_combs.and_mask_type = mask_type_normal;
            shift_combs.or_mask_type  = mask_type_none;
        }
        case riscv_shift_op_right_logical_zeros:   {
            shift_combs.and_mask_type = mask_type_invert;
            shift_combs.or_mask_type  = mask_type_none;
        }
        case riscv_shift_op_right_arithmetic:   {
            shift_combs.and_mask_type = mask_type_invert;
            shift_combs.or_mask_type  = rs1[31] ? mask_type_normal : mask_type_none;
        }
        case riscv_shift_op_left_logical_ones:   {
            if (rv_cfg_i32_bitmap_enhanced_shift_enable) {
                shift_combs.and_mask_type = mask_type_normal;
                shift_combs.or_mask_type  = mask_type_invert;
            }
        }
        case riscv_shift_op_right_logical_ones:   {
            if (rv_cfg_i32_bitmap_enhanced_shift_enable) {
                shift_combs.and_mask_type = mask_type_invert;
                shift_combs.or_mask_type  = mask_type_normal;
            }
        }
        case riscv_shift_op_left_rotate, riscv_shift_op_right_rotate, riscv_shift_op_reverse: {
            if (rv_cfg_i32_bitmap_enhanced_shift_enable) {
                shift_combs.and_mask_type = mask_type_none;
                shift_combs.or_mask_type  = mask_type_none;
            }
        }
        case riscv_shift_op_bit_insert:   {
            if (rv_cfg_i32_bitmap_enhanced_shift_enable) {
                shift_combs.and_mask_type = mask_type_normal;
                shift_combs.bb_mask_type  = bb_mask_type_bit;
                shift_combs.or_mask_type  = mask_type_rs2;
            }
        }
        case riscv_shift_op_byte_insert:   {
            if (rv_cfg_i32_bitmap_enhanced_shift_enable) {
                shift_combs.and_mask_type = mask_type_normal;
                shift_combs.bb_mask_type  = bb_mask_type_byte;
                shift_combs.or_mask_type  = mask_type_rs2;
            }
        }
        }

        /*b Find shift operands and amount; sign-extend @rshift_operand for sra, zero-extend for srl */
        shift_combs.rotate_in = rs1;
        shift_combs.shift_control = rs2[5;0];
        if (idecode.immediate_valid) { shift_combs.shift_control = idecode.immediate_shift; }

        shift_combs.shift_amount = shift_combs.shift_control;
        // shift_left must not be set for bit/byte/halfword reverse
        if (!(idecode.shift_op & riscv_shift_op_mask_right)) {
            shift_combs.shift_amount = (~shift_combs.shift_control)+1;
        }

        // swap encodings (shift_control and action)
        // 00xx0 - 000 - no swap
        // 10xx0 - 100 - swap half-words
        // 01xx0 - 010 - swap bytes, not half-words
        // 11xx0 - 110 - swap bytes, and half-words
        // 00xx1 - 001 - swap bits in bytes
        // 10xx1 - 101 - swap half-words and bits in bytes
        // 01xx1 - 011 - swap bits in bytes and bytes, not half-words
        // 11xx1 - 111 - swap bits in bytes and bytes, and half-words
        
        // half-word swap of byte swap 
        shift_combs.mask_in   = bundle(32hffffffff, 32b0);
        shift_combs.rotate_by_16 = shift_combs.rotate_in;
        if (shift_combs.shift_amount[4]) {shift_combs.rotate_by_16 = bundle(shift_combs.rotate_in[16;0], shift_combs.rotate_in[16;16]);}
        shift_combs.rotate_byte_reverse = shift_combs.rotate_by_16;
        if (shift_combs.shift_amount[3]) {
            shift_combs.rotate_byte_reverse = bundle(shift_combs.rotate_by_16[8;16], shift_combs.rotate_by_16[8;24],
                                                     shift_combs.rotate_by_16[8; 0], shift_combs.rotate_by_16[8; 8]);
        }
        shift_combs.rotate_bit_reverse = shift_combs.rotate_byte_reverse;
        if (shift_combs.shift_amount[0]) {
            for (i; 4) {
                shift_combs.rotate_bit_reverse[8;(8*i)] = bundle(shift_combs.rotate_byte_reverse[8*i+0],
                                                                 shift_combs.rotate_byte_reverse[8*i+1],
                                                                 shift_combs.rotate_byte_reverse[8*i+2],
                                                                 shift_combs.rotate_byte_reverse[8*i+3],
                                                                 shift_combs.rotate_byte_reverse[8*i+4],
                                                                 shift_combs.rotate_byte_reverse[8*i+5],
                                                                 shift_combs.rotate_byte_reverse[8*i+6],
                                                                 shift_combs.rotate_byte_reverse[8*i+7]);
            }
        }
        
        shift_combs.rotate_out = bundle(shift_combs.rotate_by_16[16;0], shift_combs.rotate_by_16) >> shift_combs.shift_amount[4;0];
        shift_combs.mask_out   = shift_combs.mask_in   >> shift_combs.shift_amount;

        /*b Determine AND and OR masks */
        shift_combs.shift_and_mask = shift_combs.mask_out[32;0];
        part_switch (shift_combs.and_mask_type) {
        case mask_type_none:   { shift_combs.shift_and_mask = -1; }
        case mask_type_invert: { shift_combs.shift_and_mask = ~shift_combs.shift_and_mask; }
        }
        if (shift_combs.shift_control==0) {
            shift_combs.shift_and_mask = -1;
        }
        if (rv_cfg_i32_bitmap_enhanced_shift_enable) {
            part_switch (shift_combs.bb_mask_type) {
            case bb_mask_type_byte: { shift_combs.shift_and_mask = shift_combs.shift_and_mask &~ (shift_combs.shift_and_mask<<8); }
            case bb_mask_type_bit:  { shift_combs.shift_and_mask = shift_combs.shift_and_mask &~ (shift_combs.shift_and_mask<<1); }
            }
        }
        shift_combs.shift_or_mask  = shift_combs.mask_out[32;0];
        if (shift_combs.shift_control==0) {
            shift_combs.shift_or_mask = 0;
        }
        part_switch (shift_combs.or_mask_type) {
        case mask_type_none:   { shift_combs.shift_or_mask = 0; }
        case mask_type_invert: { shift_combs.shift_or_mask = ~shift_combs.shift_and_mask; } // only for sllo
        case mask_type_rs2:    { shift_combs.shift_or_mask = rs2 & ~shift_combs.shift_and_mask; }
        }

        shift_combs.shift_result = (shift_combs.rotate_out[32;0] & shift_combs.shift_and_mask) | shift_combs.shift_or_mask;
        if (rv_cfg_i32_bitmap_enhanced_shift_enable) {
            if (idecode.shift_op==riscv_shift_op_reverse) {
                shift_combs.shift_result = shift_combs.rotate_bit_reverse;
            }
        }
    }

    /*b ALU operation */
    alu_operation """
    """ : {

        /*b Determine rs2 or immediate, and ditto for CSR write accesses */
        alu_combs.imm_or_rs2 = rs2;
        if (idecode.immediate_valid) { alu_combs.imm_or_rs2 = idecode.immediate; }
        alu_combs.imm_or_rs1 = rs1;
        if (idecode.immediate_valid) { alu_combs.imm_or_rs1 = idecode.immediate; }

        /*b Arithmetic operation - add with carry of rs1 with rs2+0, ~rs2+1, or imm+0, ~imm+1; used for branches and ALU op */
        alu_combs.arith_in_0 = rs1;
        alu_combs.arith_in_1 = alu_combs.imm_or_rs2;
        alu_combs.arith_carry_in = 0;
        if ((idecode.subop == riscv_subop_sub) |
            (idecode.subop == riscv_subop_slt) |
            (idecode.subop == riscv_subop_sltu)) {
            alu_combs.arith_in_1     = ~alu_combs.imm_or_rs2;
            alu_combs.arith_carry_in = 1;
        }
        if (idecode.op == riscv_op_branch) {
            alu_combs.arith_in_1     = ~rs2;
            alu_combs.arith_carry_in = 1;
        }
        if ((idecode.op == riscv_op_jalr) ||
            (idecode.op == riscv_op_mem)) {
            alu_combs.arith_in_1     = idecode.immediate;
            alu_combs.arith_carry_in = 0;
        }
        //alu_combs.arith_result      = ( bundle(1b0,alu_combs.arith_in_0) + 
        //                                bundle(1b0,alu_combs.arith_in_1) + 
        //                                bundle(32b0,alu_combs.arith_carry_in) );
        alu_combs.arith_result_32  = ( bundle(1b0,alu_combs.arith_in_0[31;0]) + 
                                        bundle(1b0,alu_combs.arith_in_1[31;0]) + 
                                        bundle(31b0,alu_combs.arith_carry_in) );
        alu_combs.carry_in_to_31 = alu_combs.arith_result_32[31];
        alu_combs.arith_result[31;0] = alu_combs.arith_result_32[31;0];
        alu_combs.arith_result[2;31] = ( bundle(1b0,alu_combs.arith_in_0[31]) + 
                                         bundle(1b0,alu_combs.arith_in_1[31]) + 
                                         bundle(1b0,alu_combs.carry_in_to_31) );
        alu_combs.arith_eq          = (alu_combs.arith_result[32;0] == 0);
        alu_combs.arith_unsigned_ge = alu_combs.arith_result[32];
        alu_combs.arith_signed_ge   = (alu_combs.carry_in_to_31 ^ alu_combs.arith_result[32])==alu_combs.arith_result[31];

        /*b Determine branch condition met */
        alu_result.branch_condition_met = 0;
        part_switch (idecode.subop) {
        case riscv_subop_beq:  {alu_result.branch_condition_met = alu_combs.arith_eq;}
        case riscv_subop_bne:  {alu_result.branch_condition_met = !alu_combs.arith_eq;}
        case riscv_subop_bgeu: {alu_result.branch_condition_met = alu_combs.arith_unsigned_ge;}
        case riscv_subop_bltu: {alu_result.branch_condition_met = !alu_combs.arith_unsigned_ge;}
        case riscv_subop_bge:  {alu_result.branch_condition_met = alu_combs.arith_signed_ge;}
        case riscv_subop_blt:  {alu_result.branch_condition_met = !alu_combs.arith_signed_ge;}
        }

        /*b Determine branch condition met */
        alu_combs.pc_plus_4    = pc + 4;
        alu_combs.pc_plus_2    = pc + 2;
        alu_combs.pc_plus_inst = idecode.is_compressed ? alu_combs.pc_plus_2 : alu_combs.pc_plus_4;
        alu_combs.pc_plus_imm = pc + idecode.immediate;
        alu_result.arith_result = alu_combs.arith_result[32;0];
        alu_result.result       = alu_combs.arith_result[32;0];
        part_switch (idecode.subop) {
        case riscv_subop_add:   { alu_result.result = alu_combs.arith_result[32;0]; }
        case riscv_subop_sub:   { alu_result.result = alu_combs.arith_result[32;0]; }
        case riscv_subop_slt:   { alu_result.result = alu_combs.arith_signed_ge   ? 0:1; }
        case riscv_subop_sltu:  { alu_result.result = alu_combs.arith_unsigned_ge ? 0:1; }
        case riscv_subop_xor:   { alu_result.result = rs1 ^ alu_combs.imm_or_rs2;}
        case riscv_subop_or:    { alu_result.result = rs1 | alu_combs.imm_or_rs2;}
        case riscv_subop_and:   { alu_result.result = rs1 & alu_combs.imm_or_rs2;}
        case riscv_subop_sll:   { alu_result.result = shift_combs.shift_result[32;0];}
        case riscv_subop_srla:  { alu_result.result = shift_combs.shift_result[32;0];}
        }
        part_switch (idecode.op) {
        case riscv_op_lui:      { alu_result.result = idecode.immediate;}
        case riscv_op_auipc:    { alu_result.result = alu_combs.pc_plus_imm;}
        case riscv_op_jal:      { alu_result.result = alu_combs.pc_plus_inst; } // jal  stores pc+2/4 ready for return in register
        case riscv_op_jalr:     { alu_result.result = alu_combs.pc_plus_inst; } // jalr stores pc+2/4 ready for return in register
        }
        alu_result.branch_target = alu_combs.pc_plus_imm;
        part_switch (idecode.op) {
        case riscv_op_jalr:     { alu_result.branch_target = bundle(alu_combs.arith_result[31;1],1b0); }
        }

        /*b CSR access write data*/
        alu_result.csr_access            = idecode.csr_access;
        alu_result.csr_access.write_data = alu_combs.imm_or_rs1;

        /*b All done */
    }

    /*b All done */
}
