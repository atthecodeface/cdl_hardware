/** Copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *   http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * @file  tb_framebuffer_teletext.cdl
 * @brief Testbench for teletext framebuffer module
 *
 * This is a simple testbench for the teletext decoder.
 */
/*a Includes */
include "srams.h"
include "teletext.h"
include "framebuffer.h"

/*a External modules */
extern module se_test_harness( clock clk "Clock for CSR reads/writes",
                               input bit reset_n,
                               output t_sram_access_req display_sram_write,
                               input t_video_bus video_bus,
                               output t_csr_request csr_request,
                               input t_csr_response csr_response
    )
{
    timing from rising clock clk   display_sram_write;
    timing from rising clock clk    csr_request;
    timing to   rising clock clk    csr_response;
    timing to   rising clock clk  video_bus;
}


/*a Module */
module tb_framebuffer_teletext( clock clk,
                                input bit reset_n
)
{

    /*b Nets */
    net t_sram_access_req display_sram_write;
    net t_video_bus video_bus;
    net t_csr_request csr_request;
    net t_csr_response csr_response;

    /*b Instantiations */
    instantiations: {
        se_test_harness th( clk <- clk,
                            display_sram_write => display_sram_write,
                            video_bus <= video_bus,
                            csr_request => csr_request,
                            csr_response <= csr_response
            );
        
        framebuffer_teletext fb( csr_clk <- clk,
                                sram_clk <- clk,
                                video_clk <- clk,
                                reset_n <= reset_n,
                                display_sram_write <= display_sram_write,
                                video_bus => video_bus,
                                csr_select_in <= 0, // uses 2 selects, from the default
                                csr_request <= csr_request,
                                csr_response => csr_response
            );
    }

    /*b All done */
}
