/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   apb_target_dprintf.cdl
 * @brief  Simple target for an APB bus to drive the dprintf request
 *
 * CDL implementation of a simple APB target to drive a dprintf request
 *
 */
/*a Includes
 */
include "dprintf.h"
include "apb.h"

/*a Types */
/*t t_apb_address
 *
 * APB address map, used to decode paddr
 */
typedef enum [2] {
    apb_address_address         = 0  "Address of register to present as the dprintf request's address",
    apb_address_data            = 1 "Eight data registers, used as the data for the dprintf request",// actually 8 to 15
    apb_address_address_commit  = 2 "Alias of the address register, with the side effect on writes of invoking the dprintf request",// actually 16 to 23
    apb_address_data_commit     = 3 "Alias of the data reigsters, with the side effect on writes of invoking the dprintf request", // actually 24 to 31
} t_apb_address;

/*t t_access
 *
 * APB access that is in progress; a decode of psel and paddr
 */
typedef enum [3] {
    access_none                  "No APB access",
    access_write_address         "Write to address register",
    access_write_address_commit  "Write to address register with a commit to invoke the dprintf request",
    access_read_address          "Read the address register",
    access_write_data            "Write a data register (selected by paddr[3;0])",
    access_write_data_commit     "Write a data register (selected by paddr[3;0]) with a commit to invoke the dprintf request",
} t_access;

/*a Module */
module apb_target_dprintf( clock clk         "System clock",
                           input bit reset_n "Active low reset",

                           input  t_apb_request  apb_request  "APB request",
                           output t_apb_response apb_response "APB response",

                           output t_dprintf_req_4 dprintf_req,
                           input  bit             dprintf_ack
    )
"""
Simple Dprintf requester with an APB interface.

A dprintf request is an address and, in this case (a @a
t_dprintf_req_4) four 64-bit data words. This is mapped to eight
32-bit data words, with data register 0 mapping to the most
significant word of the @a dprintf_req data 0 (so that data register 0
corresponds to the first text displayed as part of the dprintf).

The module provides an address register, which is the address
presented in the dprintf request. Usually for a dprintf to a teletext
framebuffer, for example, this is the address of the first character
of the output within the framebuffer.

The normal operation is to write a number of data registers, starting
with register 0, and then to write to the address register *with
commit* to invoke the dprintf.

Another method could be to have the address and bulk of the data set
up, and then a single write to a *data with commit* to, for example,
fill out a 32-bit hex value for display, invoking the dprintf (for
example if a dprintf were set up to display 'latest pc %08x', the pc
value can be written to the correct data register with commit).

The address register can be read back, in which case it has some status also:

Bits     | Meaning
---------|---------
31       | dprintf_req valid (i.e. has not been completed by dprintf slave)
15;16    | zero
16;0     | address for dprintf request.

The top bit of this register is set by a commit and cleared when the
dprintf slave acknowledges the dprintf request.

For more details on dprintf requests themselves, see the documentation in utils/src/dprintf

"""
{
    /*b Clock and reset */
    default clock clk;
    default reset active_low reset_n;

    /*b Decode APB interface */
    clocked t_access access=access_none   "Access being performed by APB";

    /*b Dprintf state */
    clocked t_dprintf_req_4 dprintf_req={*=0};

    /*b APB interface */
    apb_interface_logic """
    The APB interface is decoded to @a access when @p psel is asserted
    and @p penable is deasserted - this is the first cycle of an APB
    access. This permits the access type to be registered, so that the
    APB @p prdata can be driven from registers, and so that writes
    will occur correctly when @p penable is asserted.

    The APB read data @p prdata can then be generated based on @a
    access.
    """ : {
        /*b Decode access */
        access <= access_none;
        part_switch (apb_request.paddr[2;3]) {
        case apb_address_address: {
            access <= apb_request.pwrite ? access_write_address : access_read_address;
        }
        case apb_address_address_commit: {
            access <= apb_request.pwrite ? access_write_address_commit : access_read_address;
        }
        case apb_address_data: {
            access <= apb_request.pwrite ? access_write_data : access_none;
        }
        case apb_address_data_commit: {
            access <= apb_request.pwrite ? access_write_data_commit : access_none;
        }
        }
        if (!apb_request.psel || apb_request.penable) {
            access <= access_none;
        }

        /*b Handle APB read data */
        apb_response = {*=0, pready=1};
        part_switch (access) {
        case access_read_address: {
            apb_response.prdata = bundle(dprintf_req.valid,15b0,dprintf_req.address);
        }
        }

        /*b All done */
    }

    /*b Handle the dprintf */
    dprintf_req_logic """
    The @a dprintf_req is invalidated on an ack; it is written to by an access,
    with a commit forcing valid to 1.

    This logic is really just a set of writable registers.
    """: {
        if (dprintf_ack) {
            dprintf_req.valid <= 0;
        }
        if ((access == access_write_address_commit) || (access == access_write_data_commit)) {
            dprintf_req.valid <= 1;
        }
        if ((access == access_write_address) || (access == access_write_address_commit)) {
            dprintf_req.address <= apb_request.pwdata[16;0];
        }
        if ((access == access_write_data) || (access == access_write_data_commit)) {
            full_switch (apb_request.paddr[3;0]) {
            case 0 : {
                dprintf_req.data_0[32;32] <= apb_request.pwdata;
            }
            case 1 : {
                dprintf_req.data_0[32; 0] <= apb_request.pwdata;
            }
            case 2 : {
                dprintf_req.data_1[32;32] <= apb_request.pwdata;
            }
            case 3 : {
                dprintf_req.data_1[32; 0] <= apb_request.pwdata;
            }
            case 4 : {
                dprintf_req.data_2[32;32] <= apb_request.pwdata;
            }
            case 5 : {
                dprintf_req.data_2[32; 0] <= apb_request.pwdata;
            }
            case 6 : {
                dprintf_req.data_3[32;32] <= apb_request.pwdata;
            }
            case 7 : {
                dprintf_req.data_3[32; 0] <= apb_request.pwdata;
            }
            }
        }
    }

    /*b Done
     */
}

/*a Editor preferences and notes
mode: c ***
c-basic-offset: 4 ***
c-default-style: (quote ((c-mode . "k&r") (c++-mode . "k&r"))) ***
outline-regexp: "/\\\*a\\\|[\t ]*\/\\\*[b-z][\t ]" ***
*/
