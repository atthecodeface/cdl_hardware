/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file  teletext.cdl
 * @brief CDL implementation of a teletext decoder
 *
 * This is an implementaion of the core of a teletext decoder, for
 * arbitrary sized teletext output displays.
 *
 * The output is supplied at 12 pixels per clock (one character width)
 * The input is a byte of per clock of character data.
 *
 * The implementation does not currently support double width or
 * double size characters.
 *
 */
/*a Includes */
include "types/teletext.h"

/*a Constants */
constant integer flashing_on_count=10;
constant integer max_flashing_count=40;

/*a Types */
/*t t_color
 *
 * Three-bit color, one bit for R, G and B; this suffices for teletext
 * output
 */
typedef bit[3] t_color; // Red in [0], green in [1], blue in [2]

/*t t_character_state
 *
 * State of the character as the line is decoded, used in a number of places in the pipeline
 */
typedef struct {
    t_color background_color    "Color of background";
    t_color foreground_color    "Color of text and graphics";
    bit     flashing            "Asserted if the foreground  is flashing";
    bit     text_mode           "Asserted if the characters should be displayed as text, rather than 6-element graphics";
    bit     contiguous_graphics "Asserted if 6-element graphics should be smoothly connected; deasserted for separated elements";
    bit     double_height       "Asserted if the current character should be displayed double height";
    bit     hold_graphics_mode  "Asserted if the 'hold graphics' mode is engaged";
    bit     reset_held_graphics "Asserted if the character decodes to a control character that clears the held graphics data to space";
} t_character_state;

/*t t_timing_state
 *
 * State of the teletext frame / scanlines, to determine which part of
 * characters is to be displayed
 */
typedef struct {
    bit[5] scanline             "Scanline of character, 0 to 19; if interlaced output then 0 to 18 or 1 to 19, in twos";
    bit    last_scanline        "Asserted if on the last scanline of characters; scanline of 18 for even interlace, 19 otherwise";
    t_teletext_timings timings  "Timings as supplied by the client; effectively hsync, vsync, and how to interlace or not, etc";
    bit[6] flashing_counter     "Up-counter to determine the output color for flashing pixels; pixels turn on (foreground) if flashing_counter>flashing_on_count, counter maxes at max_flashing_count";
    bit    flash_on             "Asserted if flashing pixels should be foreground color; deasserted if they should be background";
    bit    scanline_displayed   "Asserted if there has been a valid character provided in the scanline";
} t_timing_state;

/*t t_teletext_state
 *
 * State of the line and character, valid one cycle after the input character
 */
typedef struct {
    t_teletext_character character            "Character being decoded to control the teletext state; this matches the character data being fetched by the ROM";
    t_character_state character_state         "State prior to any set-at effects of the current input character";
    bit row_contains_double_height            "Asserted if the row has had any double-height control characters";
    bit last_row_was_double_height_top        "Asserted if the last row had the top of any double-height control characters";
    bit[5] pixel_scanline                     "Scanline of the character for decode; for double height characters this differs from the timing_state scanline";
} t_teletext_state;

/*t t_teletext_combs
 *
 * Combinatorial decode of the teletext state, valid at the same time as the ROM data
 */
typedef struct {
    t_character_state set_at_character_state    "State of current character given current character state and teletext_state.character; incorporates set-at effects of the input character";
    t_character_state set_after_character_state "State of next character given current character state and teletext_state.character; incorporates set-at and set-after effects of the input character";
    bit[12] graphics_data                       "Scanline of contiguous/separated 6-element graphics data given teletext_state.character";
} t_teletext_combs;

/*t t_pixel_state
 *
 * State of the pixels, valid two cycles after the input character; depends on teletext_state and the character ROM output
 */
typedef struct {
    bit[10]              rom_scanline_data   "Two scanlines of the character data from the ROM";
    t_teletext_character character           "Character matching the scanlines from the ROM data, used for graphics decode; this matches the character data being fetched by the ROM";
    t_character_state    character_state     "Character state";
    bit[5]               pixel_scanline      "Scanline of the character for decode; for double height characters this differs from the timing_state scanline";
    bit[12]              graphics_data       "Decode of teletext_state.character as a graphics character, or possibly the held graphics";
    bit                  use_graphics_data   "Asserted if @a graphics_data should be used for the pixels, deasserted if the rom_scanline_data (possibly smoothed) should be used";
    bit[12]              held_graphics_data  "Last graphics data, unless reset by reset_held_graphics; used to replace control characters when in hold_graphics_mode";
} t_pixel_state;

/*t t_pixel_combs
 *
 * Decode of pixel state, for storing in the output_state
 */
typedef struct {
    bit[5] diagonal_0                 "SE Diagonal detection of ROM scanline data used in smoothing";
    bit[5] diagonal_1                 "SW Diagonal detection of ROM scanline data used in smoothing";
    bit[5] diagonal_2                 "NE Diagonal detection of ROM scanline data used in smoothing";
    bit[5] diagonal_3                 "NE Diagonal detection of ROM scanline data used in smoothing";
    bit[12] smoothed_scanline_data    "Smoothed scanline data generated from the two registered ROM scanlines depending on the actual scanline and the required smoothing";
} t_pixel_combs;

/*a Module teletext */
module teletext( clock clk                                "Character clock",
                 input bit reset_n                        "Active low reset",
                 input t_teletext_character    character  "Parallel character data in, with valid signal",
                 input t_teletext_timings      timings    "Timings for the scanline, row, etc",
                 output t_teletext_rom_access  rom_access "Teletext ROM access, registered output",
                 input bit[45]                 rom_data   "Teletext ROM data, valid in cycle after rom_access",
                 output t_teletext_pixels pixels          "Output pixels, three clock ticks delayed from valid data in"
       )
    /*b Documentation */
"""
This is an implementaion of the core of a presentation level 1.0
teletext decoder, for arbitrary sized teletext output displays.

The output is supplied at 12 pixels per clock (one character width)
The input is a byte of per clock of character data.

The implementation does not currently support double width or
double size characters - they are not presentation level 1.0 features.

Teletext characters are displayed from a 12x20 grid. The ROM
characters have two background rows, and then are displayed with 2
background pixels on the left, and then 10 pixels from the ROM The ROM
is actually 5x9, and it is doubled to 10x18.

The type of pixel doubling is controlled with the @a timings input. It
can be pure doubling, or smoothed. Some outputs may not want to use
the doubling, for which the best approach is to request only even
scanlines (in the @a timings) and to not smoothe, and then to select
alternate pixel color values from the output bus.

### Doubling

Doubling without smoothing can be achieved be true doubling of pixels

A simple smoothing can be performed for a pixel depending on its NSEW neighbors:


      |NN|
      |NN|
    WW|ab|EE
    WW|cd|EE
      |SS|
      |SS|

* a is filled if the pixel is filled itself, or if N&W

* b is filled if the pixel is filled itself, or if N&E

* c is filled if the pixel is filled itself, or if S&W

* d is filled if the pixel is filled itself, or if S&E

Hence one would get:

    |..|**|**|**|..|
    |..|**|**|**|..|
    |---------------
    |**|..|..|**|**|
    |**|..|..|**|**|
    |---------------
    |..|**|..|..|**|
    |..|**|..|..|**|

smoothed to:

    |..|**|**|**|..|
    |.*|**|**|**|*.|
    |---------------
    |**|*.|.*|**|**|
    |**|*.|..|**|**|
    |---------------
    |.*|**|..|.*|**|
    |..|**|..|..|**|

Or, without intervening lines:

    |..******..|
    |..******..|
    |**....****|
    |**....****|
    |..**....**|
    |..**....**|

smoothed to:

    |..******..|
    |.********.|
    |***..*****|
    |***...****|
    |.***...***|
    |..**....**|

So for even scanlines ('a' and 'b') the smoother needs row n and row n-1.

* a is set if n[x] or n[x-left]&(n-1)[x]

* b is set if n[x] or n[x-right]&(n-1)[x]

For odd scanlines ('c' and 'd') the smoother needs row n and row n+1.

* c is set if n[x] or n[x-left]&(n+1)[x]

* d is set if n[x] or n[x-right]&(n+1)[x]

This method has the unfortunate impact of smoothing two crossing lines, such as a plus:

    |....**....|     |....**....|
    |....**....|     |....**....|
    |....**....|     |....**....|
    |....**....|     |...****...|
    |**********|     |**********|
    |**********|     |**********|
    |....**....|     |...****...|
    |....**....|     |....**....|
    |....**....|     |....**....|
    |....**....|     |....**....|


Hence a better smoothing can be performed for a pixel depending on all its neighbors:

    |NW|NN|NE|
    |  |NN|  |
    |WW|ab|EE|
    |WW|cd|EE|
    |  |SS|  |
    |SW|SS|SE|

* a is filled if the pixel is filled itself, or if (N&W) but not NW

* b is filled if the pixel is filled itself, or if (N&E) but not NE

* c is filled if the pixel is filled itself, or if (S&W) but not SW

* d is filled if the pixel is filled itself, or if (S&E) but not SE

Hence one would get:

    |..|**|**|**|..|
    |..|**|**|**|..|
    |---------------
    |**|..|..|**|**|
    |**|..|..|**|**|
    |---------------
    |..|**|..|..|**|
    |..|**|..|..|**|

smoothed to:

    |..|**|**|**|..|
    |.*|**|**|**|..|
    |---------------
    |**|*.|..|**|**|
    |**|*.|..|**|**|
    |---------------
    |.*|**|..|..|**|
    |..|**|..|..|**|

Or, without intervening lines:

    |..******..|
    |..******..|
    |**....****|
    |**....****|
    |..**....**|
    |..**....**|

smoothed to:

    |..******..|
    |.*******..|
    |***...****|
    |***...****|
    |.***....**|
    |..**....**|

So for even scanlines ('a' and 'b') the smoother needs row n and row n-1.

*a is set if n[x] or (n[x-left]&(n-1)[x]) &~ (n-1)[x-left]

*b is set if n[x] or (n[x-right]&(n-1)[x]) &~ (n-1)[x-right]

For odd scanlines ('c' and 'd') the smoother needs row n and row n+1.

*c is set if n[x] or (n[x-left]&(n+1)[x]) &~ (n+1)[x-left]

*d is set if n[x] or (n[x-right]&(n+1)[x]) &~ (n+1)[x-left]


## Graphics
Graphics characters are 6 blobs on a 6x10 grid (contiguous, separated):

    |000111| |.00.11|
    |000111| |.00.11|
    |000111| |......|
    |222333| |.22.33|
    |222333| |.22.33|
    |222333| |.22.33|
    |222333| |......|
    |444555| |.44.55|
    |444555| |.44.55|
    |444555| |......|

"""
{
    /*b Defaults */
    default reset active_low reset_n;
    default clock clk;
    clocked t_timing_state    timing_state = {*=0}        "Record of which scanline and flashing, and so on; valid throughout a scanline";
    clocked t_teletext_character character_buffer = {*=0} "Character buffer to hold data while presenting ROM access";
    clocked t_teletext_state  teletext_state = {*=0}      "Teletext character state and graphics decode, one cycle later than @a character_buffer";
    comb    t_teletext_combs  teletext_combs              "Decode of the teletext state - determines graphics mode, colors, etc, and graphics character scanline data";
    clocked t_pixel_state     pixel_state={*=0}           "State from which the pixels are generated; registered data from the @a teletext_combs";
    comb    t_pixel_combs     pixel_combs                 "Decode of @a pixel_state to generate output pixels";

    /*b Timing control and character buffer stage */
    scanline_and_loading """
    First stage of the teletext pipeline.

    The character ROM controls are driven from a registered version of
    the input character. The ROM is therefore read while the
    @a teletext_combs are being evaluated, and the ROM data can be stored
    and be valid with the @a pixel_state.

    The timing logic maintains a @a scanline register, which is which
    of the twenty scanlines of the teletext character is to be
    presented. It also maintains a flashing count, which indicates
    whether flashing pixels should be foreground or background color.

    The scanline is always even for an even scanlines display - used
    for even fields of an interlaced display; for odd scanlines
    display, used in the odd fields of an interlace display, the
    scanline will always be odd. For non-interlaced displays the
    scanline increments by 1.

    If no characters are displayed on a scanline then the scanline
    counter is not updated - hence on the blank lines from the start
    of a field to the start of text, the scanline does not change, and
    so the first character row will be displayed correctly with the
    top scanline.
    """: {
        /*b Store ROM access */
        character_buffer.valid <= 0;
        if (character.valid) {
            character_buffer <= character;
        }
        rom_access = {select = character_buffer.valid,
                      address = character_buffer.character };

        /*b Record timings and update scanline */
        timing_state.timings <= timings;
        timing_state.scanline <= timing_state.scanline+2;
        if (timing_state.timings.interpolate_vertical == tvi_all_scanlines) {
            timing_state.scanline <= timing_state.scanline+1;
        }
        if (timing_state.last_scanline || timings.first_scanline_of_row) {
            timing_state.scanline <= 0;
        }
        timing_state.last_scanline <= 0;
        if (timing_state.scanline==19) {
            timing_state.last_scanline <= 1;
        }
        if ((timing_state.scanline==18) && (timing_state.timings.interpolate_vertical == tvi_even_scanlines)){
            timing_state.last_scanline <= 1;
        }

        if (!timings.first_scanline_of_row && !timings.end_of_scanline) {
            timing_state.scanline <= timing_state.scanline;
        }
        if (!timing_state.scanline_displayed) {
            timing_state.scanline <= timing_state.scanline;
        }
        if (timing_state.timings.interpolate_vertical == tvi_odd_scanlines) {
            timing_state.scanline[0] <= 1;
        }
        if (timing_state.timings.interpolate_vertical == tvi_even_scanlines) {
            timing_state.scanline[0] <= 0;
        }

        /*b Remember if anything is displayed on the scanline */
        if (timings.end_of_scanline) {
            timing_state.scanline_displayed <= 0;
        }
        if (teletext_state.character.valid) {
            timing_state.scanline_displayed <= 1;
        }

        /*b Handle a frame/field restart */
        if (timings.restart_frame) {
            timing_state.scanline_displayed <= 0;
            timing_state.scanline <= 0;
            timing_state.flashing_counter <= timing_state.flashing_counter+1;
            if (timing_state.flashing_counter==flashing_on_count) {
                timing_state.flash_on <= 1;
            }
            if (timing_state.flashing_counter==max_flashing_count) {
                timing_state.flashing_counter <= 0;
                timing_state.flash_on <= 0;
            }
        }

        /*b All done */
    }

    /*b Teletext state logic - lines up with ROM access input registers */
    teletext_state_logic """
    State at the end of the second stage of the teletext pipeline.

    Determine the scanline of the character to display, and maintain
    the teletext state for the characters as the row is analyzed.
    """: {
        /*b Store the character presented */
        teletext_state.character.valid <= 0;
        if (character_buffer.valid) {
            teletext_state.character <= character_buffer;
        }

        /*b Determine scanline - using double height if necessary */
        teletext_state.pixel_scanline <= timing_state.scanline;
        if (teletext_state.character_state.double_height) { // could use the set-at or set-after?
            teletext_state.pixel_scanline <= bundle(1b0,timing_state.scanline[4;1]);
            if (teletext_state.last_row_was_double_height_top) {
                teletext_state.pixel_scanline <= bundle(1b0,timing_state.scanline[4;1]) + 10;
            }
        }

        /*b Handle change of control state at end of character */
        if (teletext_state.character.valid) {
            teletext_state.character_state  <= teletext_combs.set_after_character_state;
            if (teletext_combs.set_at_character_state.double_height) {
                teletext_state.row_contains_double_height <= 1;
            }
        }

        /*b Handle reset of control state at end of scanline */
        if (timing_state.timings.end_of_scanline) {
            teletext_state.character_state.background_color <= 0;
            teletext_state.character_state.foreground_color <= 3b111;
            teletext_state.character_state.flashing <= 0;
            teletext_state.character_state.double_height <= 0;
            teletext_state.character_state.text_mode <= 1;
            teletext_state.character_state.hold_graphics_mode <= 0;
            teletext_state.character_state.contiguous_graphics <= 1;
        }

        /*b Handle reset of control state at end of character row */
        if (timing_state.timings.end_of_scanline && timing_state.last_scanline) {
            teletext_state.last_row_was_double_height_top <= teletext_state.row_contains_double_height ^ teletext_state.last_row_was_double_height_top;
            teletext_state.row_contains_double_height <= 0;
        }

        /*b Handle reset of control state at end of field */
        if (timing_state.timings.restart_frame) {
            teletext_state.last_row_was_double_height_top <= 0;
            teletext_state.row_contains_double_height <= 0;
        }

        /*b All done */
    }

    /*b Teletext control decode and graphics data generation during ROM access */
    teletext_control_decode """
    This is the hard work between the state at the end of stage 2 of
    the pipeline (@a teletext_state) and the end of stage 3 of the
    pipeline (@a pixel_state).

    The logic decodes the teletext state to determine the next
    teletext character state; the 'set-at' teletext info is stored in
    @a pixel_state, the 'set-after' is stored back in @a
    teletext_state.  Set-at is the notion that, for example, a 'stop
    flashing' code effects the pixels displayed for that code (it is
    set-at). Set-after is the notion that, for example, a 'red text'
    code only effects the following characters (as being in text mode,
    foreground color red).

    The graphics data that a character represents is also created;
    this will only be used if a graphics character is to be presented,
    but its generation parallels the ROM reading of the character
    scanline data so they are valid at the same time.
    
    This work is performed while the ROM data (for text characters) is
    being read.
    """: {
        /*b Decode current character while reading its contents from ROM
          note that steady, normal size, conceal, contiguous, separated, black background, new background, hold are 'set-at'
          rest are 'set-after'.
          'set-at' means it takes immediate effect for this character, 'set-after' just for the following characters
         */
        teletext_combs.set_after_character_state    = teletext_state.character_state;
        teletext_combs.set_at_character_state       = teletext_state.character_state;
        teletext_combs.set_at_character_state.reset_held_graphics = 0;
        teletext_combs.set_after_character_state.reset_held_graphics = 0; // should always be clear, only 'current' is used
        part_switch (teletext_state.character.character) {
        case 0: { // probably also the other un-interpreted <32 characters...
            teletext_combs.set_at_character_state.reset_held_graphics = 0;
        }
        case 1,2,3,4,5,6,7: {
            teletext_combs.set_after_character_state.foreground_color = teletext_state.character.character[3;0];
            teletext_combs.set_after_character_state.text_mode = 1;
            teletext_combs.set_after_character_state.hold_graphics_mode = 0; // Leaving graphics set-after, immediately... hence no hold for this
            teletext_combs.set_at_character_state.hold_graphics_mode = 0; // Although documented as set-after, it appears that the text-mode side is set-at
            teletext_combs.set_at_character_state.reset_held_graphics = !teletext_state.character_state.text_mode;
        }
        case 8: { teletext_combs.set_after_character_state.flashing = 1; }
        case 9: { // steady is set-at
            teletext_combs.set_at_character_state.flashing = 0;
            teletext_combs.set_after_character_state.flashing = 0;
        }
        case 17,18,19,20,21,22,23: {
            teletext_combs.set_after_character_state.foreground_color = teletext_state.character.character[3;0];
            teletext_combs.set_after_character_state.text_mode = 0;
            teletext_combs.set_at_character_state.reset_held_graphics = teletext_state.character_state.text_mode;
        }
        case 12: { // normal size is set-at
            teletext_combs.set_at_character_state.double_height = 0;
            teletext_combs.set_after_character_state.double_height    = 0;
            teletext_combs.set_at_character_state.reset_held_graphics = 1;
        }
        case 13: { // double height is set-after
            teletext_combs.set_at_character_state.reset_held_graphics = 1;
            teletext_combs.set_after_character_state.double_height = 1;
        }
        case 25: { // contiguous graphics is set-at
            teletext_combs.set_at_character_state.contiguous_graphics = 1;
            teletext_combs.set_after_character_state.contiguous_graphics = 1;
        }
        case 26: { // separated graphics is set-at
            teletext_combs.set_at_character_state.contiguous_graphics = 0;
            teletext_combs.set_after_character_state.contiguous_graphics = 0;
        }
        case 28: { // black background is set-at
            teletext_combs.set_at_character_state.background_color = 0;
            teletext_combs.set_after_character_state.background_color = 0;
        }
        case 29: { // new background is set-at
            teletext_combs.set_at_character_state.background_color = teletext_state.character_state.foreground_color;
            teletext_combs.set_after_character_state.background_color    = teletext_state.character_state.foreground_color;
        }
        case 30: { // hold mode is set-at
            teletext_combs.set_at_character_state.hold_graphics_mode = 1; // note that a held character is the last graphics character INCLUDING separated or not
            teletext_combs.set_after_character_state.hold_graphics_mode = 1;
        }
        case 31: { // release graphics is set-after
            teletext_combs.set_after_character_state.hold_graphics_mode = 0;
        }
        case  10, 11, 14, 15, 16, 24, 27:{
            teletext_combs.set_at_character_state.reset_held_graphics = 0;
        }
        }
        /*b Generate graphics data */
        teletext_combs.graphics_data = 12h00;
        full_switch (teletext_state.pixel_scanline[4;1]) {
        case 0, 1, 2: {
            teletext_combs.graphics_data = (teletext_state.character.character[0]?12hfc0:12h0) | (teletext_state.character.character[1]?12h03f:12h0);
        }
        case 7,8,9: {
            teletext_combs.graphics_data = (teletext_state.character.character[4]?12hfc0:12h0) | (teletext_state.character.character[6]?12h03f:12h0);
        }
        default: {
            teletext_combs.graphics_data = (teletext_state.character.character[2]?12hfc0:12h0) | (teletext_state.character.character[3]?12h03f:12h0);
        }
        }
        if (!teletext_state.character_state.contiguous_graphics) {
            teletext_combs.graphics_data[2;10] = 2b00;
            teletext_combs.graphics_data[2; 4]  = 2b00;
            part_switch (teletext_state.pixel_scanline[4;1]) {
            case 2, 6, 9: {teletext_combs.graphics_data = 0;}
            }
        }

        /*b All done */
    }

    /*b Pixel state logic - register ROM data and decoded graphics data */
    pixel_state_logic """
    Register the required scanlines of the character ROM, and store
    the appropriate graphics data to be used (if graphics is to be
    used instead of the text scanline data).

    Also, determine which color should be used as foreground - if
    flashing and the flash counter indicates 'flash off', then the
    background color replaces the foreground color in the state.
    """: {
        /*b Select scanline of ROM data for pixel and store it */
        full_switch (teletext_state.pixel_scanline[4;1]) {
        case 0: { pixel_state.rom_scanline_data <= bundle(rom_data[5;0],5b0); }
        case 1: { pixel_state.rom_scanline_data <= rom_data[10;0]; }
        case 2: { pixel_state.rom_scanline_data <= rom_data[10;5]; }
        case 3: { pixel_state.rom_scanline_data <= rom_data[10;10]; }
        case 4: { pixel_state.rom_scanline_data <= rom_data[10;15]; }
        case 5: { pixel_state.rom_scanline_data <= rom_data[10;20]; }
        case 6: { pixel_state.rom_scanline_data <= rom_data[10;25]; }
        case 7: { pixel_state.rom_scanline_data <= rom_data[10;30]; }
        case 8: { pixel_state.rom_scanline_data <= rom_data[10;35]; }
        default: { pixel_state.rom_scanline_data <= bundle(5b0,rom_data[5;40]); } // 9, and catch-all
        }
        pixel_state.pixel_scanline <= teletext_state.pixel_scanline;

        /*b Store graphics scanline data, overriding with held graphcis data if required */
        pixel_state.graphics_data     <= teletext_combs.graphics_data;
        pixel_state.use_graphics_data <= 1;
        full_switch (teletext_state.character.character[2;5]) {
        case 2b00: { // control character
            pixel_state.use_graphics_data <= 1;
            pixel_state.graphics_data     <= 0;
            if (teletext_combs.set_at_character_state.hold_graphics_mode && !teletext_combs.set_at_character_state.reset_held_graphics) {
                pixel_state.graphics_data <= pixel_state.held_graphics_data;
            }
        }
        case 2b10: { // in graphics, non-graphics character (!)
            pixel_state.use_graphics_data <= 0;
        }
        default: {
            if (teletext_state.character_state.text_mode) { // no need to use set-at/after since it is guaranteed to not be a control character
                pixel_state.use_graphics_data <= 0;
            }
        }
        }

        /*b Maintain the 'held graphics' data - last graphics data */
        if (!teletext_state.character_state.text_mode) {
            if (teletext_state.character.character[5]) {
                pixel_state.held_graphics_data <= teletext_combs.graphics_data;
            }
        }
        if (timing_state.timings.end_of_scanline) {
            pixel_state.held_graphics_data <= 0;
        }
        if (teletext_combs.set_at_character_state.reset_held_graphics) {
            pixel_state.held_graphics_data <= 0;
        }

        pixel_state.character       <= teletext_state.character; // for the valid
        if (!teletext_state.character.valid) {
            pixel_state <= pixel_state;
            pixel_state.character.valid <= 0;
        }
        pixel_state.character_state <= teletext_combs.set_at_character_state; // for the colors
        if (!timing_state.flash_on && teletext_combs.set_at_character_state.flashing) {
            pixel_state.character_state.foreground_color <= teletext_combs.set_at_character_state.background_color;
        }

        /*b All done */
    }

    /*b Pixel combinatorials - smoothe text, select text/graphics data */
    pixel_comb_logic """
    Smoothe the register scanline data, and select either that data or
    the graphics data, as determined in the previous cycle and stored
    in @a pixel_state.
    """: {
        /*b Create 'diagonals' for the character scanlines */
        pixel_combs.diagonal_0 = pixel_state.rom_scanline_data[5;5] & bundle(pixel_state.rom_scanline_data[4;0], 1b0);
        pixel_combs.diagonal_1 = pixel_state.rom_scanline_data[5;5] & bundle(1b0,pixel_state.rom_scanline_data[4;1]);
        pixel_combs.diagonal_2 = pixel_state.rom_scanline_data[5;0] & bundle(pixel_state.rom_scanline_data[4;5], 1b0);
        pixel_combs.diagonal_3 = pixel_state.rom_scanline_data[5;0] & bundle(1b0,pixel_state.rom_scanline_data[4;6]);

        pixel_combs.diagonal_0 = pixel_combs.diagonal_0 &~ bundle(pixel_state.rom_scanline_data[4;5], 1b0);
        pixel_combs.diagonal_1 = pixel_combs.diagonal_1 &~ bundle(1b0,pixel_state.rom_scanline_data[4;6]);
        pixel_combs.diagonal_2 = pixel_combs.diagonal_2 &~ bundle(pixel_state.rom_scanline_data[4;0], 1b0);
        pixel_combs.diagonal_3 = pixel_combs.diagonal_3 &~ bundle(1b0,pixel_state.rom_scanline_data[4;1]);

        /*b Create smoothed character scanline data for pixels */
        if (!pixel_state.pixel_scanline[0]) {
            pixel_combs.smoothed_scanline_data = bundle( 2b0,
                                                         pixel_state.rom_scanline_data[4]|pixel_combs.diagonal_1[4],
                                                         pixel_state.rom_scanline_data[4]|pixel_combs.diagonal_0[4],
                                                         pixel_state.rom_scanline_data[3]|pixel_combs.diagonal_1[3],
                                                         pixel_state.rom_scanline_data[3]|pixel_combs.diagonal_0[3],
                                                         pixel_state.rom_scanline_data[2]|pixel_combs.diagonal_1[2],
                                                         pixel_state.rom_scanline_data[2]|pixel_combs.diagonal_0[2],
                                                         pixel_state.rom_scanline_data[1]|pixel_combs.diagonal_1[1],
                                                         pixel_state.rom_scanline_data[1]|pixel_combs.diagonal_0[1],
                                                         pixel_state.rom_scanline_data[0]|pixel_combs.diagonal_1[0],
                                                         pixel_state.rom_scanline_data[0]|pixel_combs.diagonal_0[0]
                );
        } else {
            pixel_combs.smoothed_scanline_data = bundle( 2b0,
                                                         pixel_state.rom_scanline_data[9]|pixel_combs.diagonal_3[4],
                                                         pixel_state.rom_scanline_data[9]|pixel_combs.diagonal_2[4],
                                                         pixel_state.rom_scanline_data[8]|pixel_combs.diagonal_3[3],
                                                         pixel_state.rom_scanline_data[8]|pixel_combs.diagonal_2[3],
                                                         pixel_state.rom_scanline_data[7]|pixel_combs.diagonal_3[2],
                                                         pixel_state.rom_scanline_data[7]|pixel_combs.diagonal_2[2],
                                                         pixel_state.rom_scanline_data[6]|pixel_combs.diagonal_3[1],
                                                         pixel_state.rom_scanline_data[6]|pixel_combs.diagonal_2[1],
                                                         pixel_state.rom_scanline_data[5]|pixel_combs.diagonal_3[0],
                                                         pixel_state.rom_scanline_data[5]|pixel_combs.diagonal_2[0]
                );
        }
        if (!timing_state.timings.smoothe) {
            pixel_combs.smoothed_scanline_data = bundle( 2b0,
                                                         pixel_state.rom_scanline_data[4],pixel_state.rom_scanline_data[4],
                                                         pixel_state.rom_scanline_data[3],pixel_state.rom_scanline_data[3],
                                                         pixel_state.rom_scanline_data[2],pixel_state.rom_scanline_data[2],
                                                         pixel_state.rom_scanline_data[1],pixel_state.rom_scanline_data[1],
                                                         pixel_state.rom_scanline_data[0],pixel_state.rom_scanline_data[0] );
        }

        /*b Select text/graphics data */
        if (pixel_state.use_graphics_data) {
            pixel_combs.smoothed_scanline_data = pixel_state.graphics_data;
        }

        /*b All done */
    }

    /*b Output pixel selection, based on pixel combinatorials */
    output_pixel_selection """
    Generate output pixels by selecting the foreground or background
    color, based on either the character data or the graphics data
    which is presented as @a pixel_combs.smoothed_scanline_data.

    For flashing colors the foreground_color should have already been
    changed (if flash off) to match the background color, so no need
    to account for flashing here.
    """: {
        /*b Generate colored pixels */
        pixels.red = 0;
        pixels.blue = 0;
        pixels.green = 0;

        for (i; 12) {
            pixels.red[i]   = pixel_state.character_state.background_color[0];
            pixels.green[i] = pixel_state.character_state.background_color[1];
            pixels.blue[i]  = pixel_state.character_state.background_color[2];
            if (pixel_combs.smoothed_scanline_data[i]) {
                pixels.red[i]   = pixel_state.character_state.foreground_color[0];
                pixels.green[i] = pixel_state.character_state.foreground_color[1];
                pixels.blue[i]  = pixel_state.character_state.foreground_color[2];
            }
        }
        pixels.valid         = pixel_state.character.valid;
        pixels.last_scanline = timing_state.last_scanline;
    }

    /*b All done */
}
