/** Copyright (C) 2019,  Gavin J Stark.  All rights reserved.
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *   http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * @file  tb_clocking.cdl
 * @brief Testbench for numerous clocking modules
 *
 */
/*a Includes */
include "types/timer.h"
include "clocking/clock_timer_modules.h"

/*a External modules */
extern module se_test_harness( clock clk,
                               output t_timer_control   master_timer_control,
                               output t_timer_control   slave_timer_control,
                               input  t_timer_value     master_timer_value,
                               input  t_timer_value     slave_timer_value,
                               input  t_timer_sec_nsec  master_timer_sec_nsec,
                               input  t_timer_sec_nsec  slave_timer_sec_nsec
    )
{
    timing from rising clock clk master_timer_control, slave_timer_control;
    timing to   rising clock clk master_timer_value, slave_timer_value, master_timer_sec_nsec, slave_timer_sec_nsec;
}

/*a Module */
module tb_clock_timer( clock clk,
                       clock slave_clk,
                       input bit reset_n
)
{

    /*b Nets */
    net t_timer_control   master_timer_control;
    net t_timer_control   slave_timer_control;
    net t_timer_control   slave_timer_control_out;
    net t_timer_value     master_timer_value;
    net t_timer_value     slave_timer_value;
    net t_timer_sec_nsec  master_timer_sec_nsec;
    net t_timer_sec_nsec  slave_timer_sec_nsec;

    /*b Instantiations */
    instantiations: {
        se_test_harness th( clk <- clk,
                            master_timer_control => master_timer_control,
                            slave_timer_control  => slave_timer_control,
                            master_timer_value   <= master_timer_value,
                            slave_timer_value    <= slave_timer_value,
                            master_timer_sec_nsec <= master_timer_sec_nsec,
                            slave_timer_sec_nsec  <= slave_timer_sec_nsec
            );
        clock_timer ckt( clk <- clk, reset_n <= reset_n,
                         timer_control <= master_timer_control,
                         timer_value   => master_timer_value
            );
        clock_timer_async ckts( master_clk <- clk, master_reset_n <= reset_n,
                                slave_clk <- slave_clk, slave_reset_n <= reset_n,
                                master_timer_control <= master_timer_control,
                                master_timer_value   <= master_timer_value,
                                slave_timer_control_in  <= slave_timer_control,
                                slave_timer_control_out => slave_timer_control_out,
                                slave_timer_value    => slave_timer_value
            );
        clock_timer_as_sec_nsec ctasn_m( clk <- clk,
                                 reset_n <= reset_n,
                                 timer_control <= master_timer_control,
                                 timer_value   <= master_timer_value,
                                 timer_sec_nsec => master_timer_sec_nsec
            );
        clock_timer_as_sec_nsec ctasn_s( clk <- slave_clk,
                                 reset_n <= reset_n,
                                 timer_control <= slave_timer_control_out,
                                 timer_value   <= slave_timer_value,
                                 timer_sec_nsec => slave_timer_sec_nsec
            );
    }

    /*b All done */
}
