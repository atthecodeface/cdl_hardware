/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   riscv_minimal.cdl
 * @brief  Minimal RISC-V implementation ported to CDL
 *
 * CDL implementation of 3-stage minimal RISC-V teaching implementation
 *
 * This is a three stage pipeline implementation (not including
 * instruction fetch itself).
 *
 * The first stage is decode and register file read
 *
 * The second stage is data forwarding, ALU, data memory request, CSR access, conditional branching, jump table branching and traps.
 *
 * The third stage is data memory read (the memory is doing stuff, the CPU is not), rotating the data read and merging (for unaligned transfers)
 *
 * The end of the third stage is register file writeback; there is a register in RFW for memory data written to last register
 *
 *
 * Decode stage: Instruction register, PC, valid
 *
 * decode i32/i32c -> rfr ports -> rf mux
 *
 * ALU stage: RFR values, decoded instruction, PC, valid, predicted_taken, cycle of instruction
 *
 * ALU result/mem result/RFR mux -> ALU operation -> Dmem access request -> jump
 *
 * Mem stage: ALU result, MEM request in progress, valid, rd, rd_valid
 *
 * Mem in progress -> data read -> rotate data
 *
 * RFW stage: MEM result, RF
 *
 */

/*a Includes
 */
include "riscv_internal_types.h"
include "riscv.h"
include "riscv_submodules.h"

/*a Constants
 */
constant integer INITIAL_PC=0x80000000;
constant integer i32c_force_disable=0;
constant integer coproc_force_disable=0;

/*a Types
 */
/*t t_ifetch_combs
 *
 * Combinatorials for the instruction fetch
 */
typedef struct {
    bit request;
    bit[32] address;
    bit sequential;
} t_ifetch_combs;

/*t t_dec_state */
typedef struct {
    bit enable                   "Asserted if execution is enabled, deasserted at reset";
    t_riscv_i32_inst instruction   "Fetched instruction, ready for decode, register fetch, execute and writeback";
    bit valid                    "Asserted if @instruction is a valid fetched instruction, whether misaligned or not";
    bit illegal_pc               "Asserted if a valid @instruction is a fetched instruction from a badly aligned PC";
    bit[32] pc                   "PC of the fetched instruction";
    bit     fetch_sequential     "Asserted if?";
} t_dec_state;

/*t t_dec_combs
 *
 * Combinatorials of the decode state
 */
typedef struct {
    t_riscv_i32_decode idecode;

    t_riscv_word   rs1;
    t_riscv_word   rs2;

    bit[32] pc_plus_4;
    bit[32] pc_plus_2;
    bit[32] pc_plus_inst;
    bit[32] pc_branch_target;
    bit predict_branch;

    bit[32] fetch_next_pc;
    bit[32] pc_if_mispredicted   "PC of the next instruction if branch prediction is incorrect";
    bit     fetch_sequential;

    bit rs1_from_alu;
    bit rs1_from_mem;
    bit rs2_from_alu;
    bit rs2_from_mem;

} t_dec_combs;

/*t t_alu_state */
typedef struct {
    bit valid;
    bit first_cycle              "Asserted if first cycle of an instruction execution (so instruction can be interrupted)";
    t_riscv_i32_decode idecode;
    bit[32] pc                   "PC of the fetched instruction";
    bit illegal_pc               "Asserted if a valid @instruction is a fetched instruction from a badly aligned PC";
    bit[32] pc_if_mispredicted   "PC of the next instruction if branch prediction is incorrect";
    bit predicted_branch         "Asserted if instruction decode predicted this is a taken branch";
    bit rs1_from_alu;
    bit rs1_from_mem;
    bit rs2_from_alu;
    bit rs2_from_mem;
    t_riscv_word   rs1;
    t_riscv_word   rs2;

    t_riscv_i32_inst debug_instruction    "Decoded instruction, for trace only";
} t_alu_state;

/*t t_alu_combs
 *
 * Combinatorials of the ALU stage
 */
typedef struct {
    bit valid_legal              "Asserted if @instruction is a valid fetched instruction on a valid alignment";
    bit blocked_by_mem           "Must qualify with valid; asserted if the ALU instruction cannot start because it uses a result of the memory stage";
    bit cannot_start             "Asserted if the instruction is blocked from starting; ignored unless valid and first_cycle; can be because of blocked_by_mem or coprocessor not ready";
    bit cannot_complete          "Asserted if the ALU has a valid instruction that either cannot be started or cannot complete";
    bit flush_pipeline;
    bit[32] next_pc;
    t_riscv_word   rs1;
    t_riscv_word   rs2;
    bit[2]  word_offset;
    bit reading;
    bit[2] read_data_rotation;
    bit[4] read_data_byte_clear;
    bit[4] read_data_byte_enable;
    bit branch_taken;
    bit trap;
    bit mret;
    bit jalr;
    t_riscv_trap_cause trap_cause;
    bit[32] trap_value;
    t_riscv_csr_access csr_access;
    t_riscv_word result_data;
    bit dmem_misaligned          "Asserted if the dmem address offset in a word does not match the size of the decoded access, whether the instruction is valid or not";
    bit dmem_multicycle          "Asserted if dmem_misaligned and it would take 2 transactions to satisfy the memory operation, whether the instruction is valid or not";
} t_alu_combs;

/*t t_mem_state */
typedef struct {
    bit valid                   "Asserted if the state here is valid";
    t_riscv_word alu_result     "Result from the last alu stage; this will be combined with memory result to be stored in RF";
    bit rd_written              "Asserted if Rd is to be written to (with result of memory or ALU)";
    bit rd_from_mem             "Asserted if Rd is to be written to with result of memory - so a following instruction must wait until this one reaches RFW";
    bit[5] rd                   "Destination register used by the instruction (if valid and rd_written are asserted)";
    bit reading                 "Asserted if the memory is reading and data should be merged with previous mem result";
    bit[4] byte_clear           "Bytes of current rfw_state.mem_result to clear in merging with memory read data for memory result (for unaligned reads)";
    bit[4] byte_enable          "Bytes of memory read data to be merged with current rfw_state.mem_result for memory result (for unaligned reads)";
    bit[2] rotation             "Number of bytes to rotate memory read data right by to get it in to correct byte alignment before merging";
    bit sign_extend_byte;
    bit sign_extend_half;
} t_mem_state;

/*t t_mem_combs
 *
 * Combinatorials of the memory stage
 */
typedef struct {
    t_riscv_word aligned_data;
    t_riscv_word memory_data;
    t_riscv_word result_data;
} t_mem_combs;

/*t t_rfw_state */
typedef struct {
    bit valid                   "Asserted if the state here is valid";
    t_riscv_word mem_result     "Result from the last mem stage; this was written to the RF (if required) at the same time it was stored here";
    bit rd_written              "Asserted if Rd of the RF was written to";
    bit[5] rd                   "Destination register used by the instruction (if valid and rd_written are asserted)";
} t_rfw_state;

/*a Module
 */
module riscv_i32c_pipeline3( clock clk,
                             input bit reset_n,
                             output t_riscv_mem_access_req  dmem_access_req,
                             input  t_riscv_mem_access_resp dmem_access_resp,
                             output t_riscv_fetch_req       ifetch_req,
                             input  t_riscv_fetch_resp      ifetch_resp,
                             output t_riscv_i32_coproc_controls  coproc_controls,
                             input t_riscv_i32_coproc_response   coproc_response,
                             input  t_riscv_config          riscv_config,
                             output t_riscv_i32_trace       trace
)
"""
This is just the processor pipeline, using thress stages for execution.

The decode and RFR is performed in the first stage

The ALU execution (and coprocessor execution) is performed in the second stage

Memory operations are performed in the third stage

Register file is written at the end of the third stage; there is a RFW stage to
forward data from RFW back to execution.

Instruction fetch
-----------------

The instruction fetch request for the next cycle is put out just after
the ALU stage logic, which may be a long time into the cycle
(althought the design keeps this to a minimum); the fetch data
response presents the instruction fetched at the end of the cycle,
where it is registered for execution.

The instruction fetch response must then be valid combinatorially
based on the instruction fetch request.

Data memory access
------------------

The data memory request is presented in the ALU stage, for an access
to complete during the memory stage.

To support simple synchronous memory operation the data memory access
includes valid write data in the same cycle as the request.

The data memory response is valid one cycle later than a request. This
includes a wait signal. The external memory subsystem, therefore, is a
two stage pipeline. The wait signal controls whether an access
completes, but not if an access can be taken (except indirectly).

Hence external logic must always either register a request or
guarantee not to assert wait.

An example implementation of could be
    dmem_access_resp.wait = fn ( access_in_progress );
    access_can_be_taken = (!access_in_progress.valid) || (!dmem_access_resp.wait);
    if (access_can_be_taken) {
      access_in_progress <= dmem_access_req;
    }
}

"""
{

    /*b State and comb
     */
    default clock clk;
    default reset active_low reset_n;

    clocked t_riscv_word[32] registers={*=-1} "Register 0 is tied to 0 - so it is written on every cycle to zero...";

    comb    t_ifetch_combs         ifetch_combs;
    net     t_riscv_i32_decode     idecode_i32;
    net     t_riscv_i32_decode     idecode_i32c;
    net     t_riscv_i32_alu_result alu_result;

    comb t_dec_combs dec_combs;
    comb t_alu_combs alu_combs;
    comb t_mem_combs mem_combs;
    clocked t_dec_state     dec_state={*=0, pc=INITIAL_PC};
    clocked t_alu_state     alu_state={*=0};
    clocked t_mem_state     mem_state={*=0};
    clocked t_rfw_state     rfw_state={*=0};
    comb t_riscv_i32_coproc_response   coproc_response_cfg "Coprocessor response masked out if configured off";

    comb t_riscv_csr_controls csr_controls;
    net t_riscv_csr_data csr_data;
    net t_riscv_csrs_minimal csrs;

    /*b Ifetch request
     */
    instruction_fetch_request
    """
    The instruction fetch request derives from the decode stage for
    conditional branches (predicted taken if backwards) and for
    unconditional branches.

    If the decode stage is invalid (i.e. it does not have a
    valid instruction to decode) then the current decode stage PC is requested.

    However, if the execute stage is valid and
    a trap is taken, or a forward conditional branch is taken or a
    backward conditional branch is not taken or a jump table branch is
    taken, then the execute stage result pc has to be used.

    This request may be for any 16-bit aligned address, and two
    successive 16-bit words from that request must be presented,
    aligned to bit 0.

    """:
    {
        ifetch_combs.address        = dec_combs.fetch_next_pc;
        ifetch_combs.sequential     = dec_combs.fetch_sequential;
        if (!dec_state.valid) {
            ifetch_combs.address    = dec_state.pc;
            ifetch_combs.sequential = dec_state.fetch_sequential;
        }

        if (alu_state.valid && alu_combs.flush_pipeline) {
            ifetch_combs.address    = alu_combs.next_pc;
            ifetch_combs.sequential = 0;
        }

        ifetch_combs.request = dec_state.enable;

        ifetch_req             = {*=0};
        ifetch_req.valid       = ifetch_combs.request;
        ifetch_req.sequential  = ifetch_combs.sequential;
        ifetch_req.address     = ifetch_combs.address;
    }

    /*b Decode, RFR stage
     */
    decode_rfr_stage """
    The decode/RFR stage decodes an instruction, follows unconditional
    branches and backward conditional branches (to generate the next
    PC as far as decode is concerned), determines register forwarding
    required, reads the register file.
    """: {
        /*b Enable operation (zeroed in reset) */
        dec_state.enable <= 1;

        /*b Instruction register - note all PC value are legal (bit 0 is cleared automatically though) */
        dec_state.valid <= 0;
        if (alu_combs.cannot_complete && dec_state.valid) {
            dec_state <= dec_state;
        } elsif (ifetch_req.valid) {
            if (ifetch_resp.valid) {
                dec_state.valid <= 1;
                dec_state.instruction <= {data=ifetch_resp.data, mode=rv_mode_machine};
                dec_state.illegal_pc <= 0;
            }
            dec_state.pc               <= ifetch_req.address;
            dec_state.fetch_sequential <= ifetch_req.sequential;
        }

        /*b Decode instruction */
        riscv_i32_decode decode_i32( instruction <= dec_state.instruction,
                                     idecode     => idecode_i32,
                                     riscv_config      <= riscv_config );

        riscv_i32c_decode decode_i32c( instruction <= dec_state.instruction,
                                       idecode      => idecode_i32c,
                                       riscv_config      <= riscv_config );

        /*b Select decode */
        dec_combs.idecode = idecode_i32;
        if ((!i32c_force_disable) && riscv_config.i32c) {
            if (dec_state.instruction.data[2;0]!=2b11) {
                dec_combs.idecode = idecode_i32c;
            }
        }

        /*b Register read */
        dec_combs.rs1 = registers[dec_combs.idecode.rs1]; // note that register 0 is ALWAYS 0 anyway
        dec_combs.rs2 = registers[dec_combs.idecode.rs2]; // note that register 0 is ALWAYS 0 anyway

        /*b Detect unconditional branches and backward conditional branches */
        dec_combs.pc_plus_4      = dec_state.pc + 4;
        dec_combs.pc_plus_2      = dec_state.pc + 2;
        dec_combs.pc_plus_inst   = dec_combs.idecode.is_compressed ? dec_combs.pc_plus_2 : dec_combs.pc_plus_4;
        dec_combs.pc_branch_target  = dec_state.pc + dec_combs.idecode.immediate;
        dec_combs.predict_branch = 0;

        part_switch (dec_combs.idecode.op) {
        case riscv_op_branch:   { dec_combs.predict_branch = dec_combs.idecode.immediate[31]; }
        case riscv_op_jal:      { dec_combs.predict_branch = 1; }
        }

        dec_combs.fetch_next_pc      = dec_combs.pc_plus_inst;
        dec_combs.fetch_sequential   = 1;
        dec_combs.pc_if_mispredicted = dec_combs.pc_branch_target;
        if (dec_combs.predict_branch) {
            dec_combs.fetch_next_pc      = dec_combs.pc_branch_target;
            dec_combs.fetch_sequential   = 0;
            dec_combs.pc_if_mispredicted = dec_combs.pc_plus_inst;
        }
        
        /*b Register forwarding determination */
        dec_combs.rs1_from_alu = 0;
        dec_combs.rs1_from_mem = 0;
        dec_combs.rs2_from_alu = 0;
        dec_combs.rs2_from_mem = 0;
        if ((mem_state.rd == dec_combs.idecode.rs1) && mem_state.rd_written) {
            dec_combs.rs1_from_mem = 1;
        }
        if ((alu_state.idecode.rd == dec_combs.idecode.rs1) && alu_state.idecode.rd_written) {
            dec_combs.rs1_from_alu = 1;
        }
        if ((mem_state.rd == dec_combs.idecode.rs2) && mem_state.rd_written) {
            dec_combs.rs2_from_mem = 1;
        }
        if ((alu_state.idecode.rd == dec_combs.idecode.rs2) && alu_state.idecode.rd_written) {
            dec_combs.rs2_from_alu = 1;
        }
    }

    /*b ALU (execute) stage registers (alu_state)
     */
    alu_stage """
    The ALU stage does data forwarding, ALU operation, conditional branches, CSR accesses, memory request
    """: {
        /*b Record state */
        alu_state.valid <= 0;
        alu_state.idecode.rd_written <= 0; // Ensure it is cleared if invalid
        if (alu_combs.cannot_complete) {
            if (!alu_combs.cannot_start) {
                alu_state.first_cycle <= 0;
            }
            alu_state <= alu_state;
            alu_state.rs1_from_alu <= 0;
            alu_state.rs2_from_alu <= 0;
            alu_state.rs1_from_mem <= alu_state.rs1_from_alu;
            alu_state.rs2_from_mem <= alu_state.rs2_from_alu;
            if (alu_state.rs1_from_mem) {
                alu_state.rs1 <= rfw_state.mem_result;
            }
            if (alu_state.rs2_from_mem) {
                alu_state.rs2 <= rfw_state.mem_result;
            }
        } elsif (dec_state.valid && !alu_combs.flush_pipeline) {
            alu_state.valid               <= 1;
            alu_state.first_cycle         <= 1;
            alu_state.illegal_pc          <= dec_state.illegal_pc;
            alu_state.idecode             <= dec_combs.idecode;
            alu_state.pc                  <= dec_state.pc;
            alu_state.pc_if_mispredicted  <= dec_combs.pc_if_mispredicted;
            alu_state.predicted_branch    <= dec_combs.predict_branch;
            alu_state.rs1                 <= dec_combs.rs1;
            alu_state.rs2                 <= dec_combs.rs2;
            alu_state.rs1_from_alu        <= dec_combs.rs1_from_alu;
            alu_state.rs1_from_mem        <= dec_combs.rs1_from_mem;
            alu_state.rs2_from_alu        <= dec_combs.rs2_from_alu;
            alu_state.rs2_from_mem        <= dec_combs.rs2_from_mem;

            alu_state.debug_instruction   <= dec_state.instruction;
        }
    }

    /*b ALU (execute) stage logic (alu_combs)
     */
    alu_stage_logic """
    The ALU stage does data forwarding, ALU operation, conditional branches, CSR accesses, memory request
    """: {
        alu_combs.valid_legal = alu_state.valid && !alu_state.idecode.illegal;

        /*b Data forwarding */
        alu_combs.rs1 = alu_state.rs1;
        alu_combs.blocked_by_mem = 0;
        if (alu_state.rs1_from_mem) {
            alu_combs.rs1 = rfw_state.mem_result;
        }
        if (alu_state.rs1_from_alu) {
            alu_combs.rs1 = mem_state.alu_result;
            if (mem_state.rd_from_mem) {
                alu_combs.blocked_by_mem = alu_state.idecode.rs1_valid;
            }
        }
        alu_combs.rs2 = alu_state.rs2;
        if (alu_state.rs2_from_mem) {
            alu_combs.rs2 = rfw_state.mem_result;
        }
        if (alu_state.rs2_from_alu) {
            alu_combs.rs2 = mem_state.alu_result;
            if (mem_state.rd_from_mem) {
                alu_combs.blocked_by_mem = alu_state.idecode.rs2_valid;
            }
        }
        alu_combs.cannot_start    = alu_combs.blocked_by_mem || coproc_response_cfg.cannot_start;
        alu_combs.cannot_complete = alu_combs.cannot_start   || coproc_response_cfg.cannot_complete;

        /*b Execute ALU stage */
        riscv_i32_alu alu( idecode <= alu_state.idecode,
                           pc  <= alu_state.pc,
                           rs1 <= alu_combs.rs1,
                           rs2 <= alu_combs.rs2,
                           alu_result => alu_result );

        /*b Minimal CSRs */
        csr_controls = {*=0};
        csr_controls.retire      = alu_combs.valid_legal;
        csr_controls.timer_inc   = 1;

        alu_combs.csr_access = alu_state.idecode.csr_access;
        if (!alu_combs.valid_legal) {
            alu_combs.csr_access.access = riscv_csr_access_none;
        }
        riscv_csrs_minimal csrs( clk <- clk,
                                 reset_n <= reset_n,
                                 csr_access     <= alu_combs.csr_access,
                                 csr_write_data <= alu_state.idecode.illegal ? bundle(27b0, alu_state.idecode.rs1) : alu_combs.rs1,
                                 csr_data       => csr_data,
                                 csr_controls   <= csr_controls,
                                 csrs => csrs);

        /*b ALU stage result */
        alu_combs.result_data = alu_result.result | coproc_response_cfg.result;
        if (coproc_response_cfg.result_valid) {
            alu_combs.result_data = coproc_response_cfg.result;
        }
        if (alu_state.idecode.csr_access.access != riscv_csr_access_none) {
            alu_combs.result_data = csr_data.read_data;
        }

        /*b Memory access handling */
        dmem_access_req.read_enable  = (alu_state.idecode.op == riscv_op_load);
        dmem_access_req.write_enable = (alu_state.idecode.op == riscv_op_store);
        if (!alu_state.valid) {
            dmem_access_req.read_enable  = 0;
            dmem_access_req.write_enable = 0;
        }
        alu_combs.reading = dmem_access_req.read_enable;

        dmem_access_req.address   = alu_result.arith_result;
        alu_combs.word_offset     = alu_result.arith_result[2;0];
        alu_combs.dmem_misaligned = (alu_combs.word_offset!=0); // valid for words
        alu_combs.dmem_multicycle = (alu_combs.word_offset!=0); // valid for words
        alu_combs.read_data_rotation = alu_combs.word_offset;
        alu_combs.read_data_byte_enable = 4hf;
        alu_combs.read_data_byte_clear  = 4hf;
        part_switch (alu_state.idecode.memory_width) {
        case mw_byte: {
            dmem_access_req.byte_enable  = 4h1 << alu_combs.word_offset;
            alu_combs.read_data_byte_enable = 4h1;
            alu_combs.dmem_misaligned = 0;
            alu_combs.dmem_multicycle = 0;
        }
        case mw_half: {
            dmem_access_req.byte_enable  = 4h3 << alu_combs.word_offset;
            alu_combs.read_data_byte_enable = 4h3;
            alu_combs.dmem_misaligned = alu_combs.word_offset[0];
            alu_combs.dmem_multicycle = (alu_combs.word_offset==2b11);
        }
        default: {
            dmem_access_req.byte_enable  = 4hf << alu_combs.word_offset;
            alu_combs.dmem_misaligned = (alu_combs.word_offset!=0);
            alu_combs.dmem_multicycle = (alu_combs.word_offset!=0);
        }
        }

        dmem_access_req.write_data = alu_combs.rs2;
        full_switch (alu_combs.word_offset) {
        case 2b00: { dmem_access_req.write_data = alu_combs.rs2; }
        case 2b01: { dmem_access_req.write_data = bundle(alu_combs.rs2[24; 0], alu_combs.rs2[ 8;24]); }
        case 2b10: { dmem_access_req.write_data = bundle(alu_combs.rs2[16; 0], alu_combs.rs2[16;16]); }
        case 2b11: { dmem_access_req.write_data = bundle(alu_combs.rs2[ 8; 0], alu_combs.rs2[24; 8]); }
        }

        /*b Determine whether to trap

          Trap sources are:

          software interrupt (ecall)
            epc <= address of instruction (even if it was a compressed inst)
          debug 
            lowest priority:  single step
            next priority:    debugger requested
            next priority:    ebreak with DCSR[ebreak*] set
              epc <= address of instruction (even if it was a compressed inst)
            highest priority: trigger with action=enter-debug-mode          
          unaligned instruction fetch
          unaligned data operation
            load or atomic/store

         */
        alu_combs.trap = 0;
        alu_combs.trap_cause = 0;
        alu_combs.trap_value = 0;
        part_switch (alu_state.idecode.op) {
        case riscv_op_system:   {
            if (alu_state.idecode.subop==riscv_subop_ecall) {
                alu_combs.trap = 1;
                alu_combs.trap_cause = riscv_trap_cause_mecall;
            }
            if (alu_state.idecode.subop==riscv_subop_ebreak) {
                alu_combs.trap = 1;
                alu_combs.trap_cause = riscv_trap_cause_breakpoint;
                alu_combs.trap_value = alu_state.pc; // WHY???
            }
        }
        }
        if (alu_state.idecode.illegal) {
            alu_combs.trap = 1;
            alu_combs.trap_cause = riscv_trap_cause_illegal_instruction;
            alu_combs.trap_value = alu_state.debug_instruction.data; // OPTIONAL???
        }
        if (alu_state.illegal_pc) {
            alu_combs.trap       = 1;
            alu_combs.trap_cause = riscv_trap_cause_instruction_misaligned;
            alu_combs.trap_value = alu_state.pc;
        }

        csr_controls.trap_cause = alu_combs.trap_cause;
        csr_controls.trap       = 0;
        csr_controls.trap_pc    = alu_state.pc;
        csr_controls.trap_value = alu_combs.trap_value;
        if (alu_combs.trap) {
            csr_controls.trap       = alu_state.valid;
        }

        /*b Determine whether branch would be taken and find next PC */
        alu_combs.branch_taken = 0;
        alu_combs.mret = 0;
        alu_combs.jalr = 0;
        part_switch (alu_state.idecode.op) {
        case riscv_op_branch:   { alu_combs.branch_taken = alu_result.branch_condition_met; }
        case riscv_op_jal:      { alu_combs.branch_taken=1; }
        case riscv_op_jalr:     {
            alu_combs.jalr = 1;
        }
        case riscv_op_system:   {
            if (alu_state.idecode.subop==riscv_subop_mret) {
                alu_combs.mret = 1;
            }
        }
        }

        alu_combs.flush_pipeline = 0;
        alu_combs.next_pc        = alu_state.pc_if_mispredicted; // only used if flushing
        if (alu_combs.branch_taken) { // branch IS to be taken - flush if a branch was not predicted
            alu_combs.flush_pipeline = !alu_state.predicted_branch;
        } else { // branch is NOT to be taken - flush if a branch was predicted
            alu_combs.flush_pipeline = alu_state.predicted_branch;
        }
        if (alu_combs.jalr) {
            alu_combs.flush_pipeline = 1;
            alu_combs.next_pc = alu_result.arith_result;
        }
        if (alu_combs.mret) { // must change mode and set interrupt enables appropriately!
            alu_combs.flush_pipeline = 1;
            alu_combs.next_pc = csrs.mepc;
        }
        if (alu_combs.trap) {
            alu_combs.flush_pipeline = 1;
            alu_combs.next_pc = csrs.mtvec;
        }
        if (!alu_state.valid || alu_combs.cannot_complete) {
            alu_combs.flush_pipeline = 0;
        }

    }

    /*b Memory stage
     */
    memory_stage """
    The memory access stage is when the memory is performing a read

    When unaligned accesses are supported this will merge two reads
    using multiple cycles

    This is a single cycle, with committed transactions only being
    valid

    If the memory is performing a read then the memory data is rotated
    and presented as the result; otherwise the ALU result is passed
    through.

    """: {
        /*b State - tie some things down so that data path does not toggle so much */
        mem_state.valid        <= 0;
        mem_state.reading      <= 0;
        mem_state.rd_written   <= 0;
        mem_state.rd_from_mem  <= 0;
        mem_state.rotation     <= 0;
        mem_state.byte_enable  <= 0;
        mem_state.byte_clear   <= 4hf;
        if (alu_combs.valid_legal && !alu_combs.cannot_complete) {
            mem_state.valid        <= 1;
            mem_state.reading      <= alu_combs.reading;
            mem_state.rotation     <= alu_combs.read_data_rotation;
            mem_state.byte_enable  <= alu_combs.read_data_byte_enable;
            mem_state.byte_clear   <= alu_combs.read_data_byte_clear;
            mem_state.rd_written   <= alu_state.idecode.rd_written;
            if (alu_combs.reading && alu_state.idecode.rd_written) {
                mem_state.rd_from_mem <= 1;
            }
            mem_state.rd           <= alu_state.idecode.rd;
            mem_state.alu_result   <= alu_combs.result_data;
            mem_state.sign_extend_half <= ((!alu_state.idecode.memory_read_unsigned) && (alu_state.idecode.memory_width== mw_half));
            mem_state.sign_extend_byte <= ((!alu_state.idecode.memory_read_unsigned) && (alu_state.idecode.memory_width== mw_byte));
        }

        /*b Memory read handling */
        mem_combs.aligned_data = dmem_access_resp.read_data;
        full_switch (mem_state.rotation) {
        case 2b00: {
            mem_combs.aligned_data = dmem_access_resp.read_data;
        }
        case 2b01: {
            mem_combs.aligned_data = bundle(dmem_access_resp.read_data[ 8;0], dmem_access_resp.read_data[24; 8]);
        }
        case 2b10: {
            mem_combs.aligned_data = bundle(dmem_access_resp.read_data[16;0], dmem_access_resp.read_data[16;16]);
        }
        case 2b11: {
            mem_combs.aligned_data = bundle(dmem_access_resp.read_data[24;0], dmem_access_resp.read_data[ 8;24]);
        }
        }
        mem_combs.memory_data = mem_combs.aligned_data;
        for (i; 4) {
            mem_combs.memory_data[8;8*i] = ( (mem_state.byte_clear[i]?8b0:mem_state.alu_result[8;8*i]) |
                                             (mem_state.byte_enable[i]?mem_combs.aligned_data[8;8*i]:8b0) );
        }
        if (mem_state.sign_extend_byte && mem_combs.memory_data[7])  { mem_combs.memory_data[24;8]  = -1; }
        if (mem_state.sign_extend_half && mem_combs.memory_data[15]) { mem_combs.memory_data[16;16] = -1; }

        /*b Memory result mux */
        mem_combs.result_data = mem_state.alu_result;
        if (mem_state.reading) {
            mem_combs.result_data = mem_combs.memory_data;
        }
    }

    /*b RFW 'stage'
     */
    rfw_stage """
    The RFW stage takes the memory read data and memory stage internal data,
    and combines them, preparing the result for the register file (written at the end of the clock)
    """: {
        /*b RFW state */
        rfw_state.valid        <= 0;
        rfw_state.rd_written   <= 0;
        if (mem_state.valid) {
            rfw_state.valid        <= 1;
            rfw_state.rd_written   <= mem_state.rd_written;
            rfw_state.rd           <= mem_state.rd;
            rfw_state.mem_result   <= mem_combs.result_data;
            if (mem_state.rd_written) {
                registers[mem_state.rd] <= mem_combs.result_data;
            }
        }
        registers[0] <= 0; // register 0 is always zero...
    }

    /*b Coprocessor interface */
    coprocessor_interface """
    Drive the coprocessor controls unless disabled; mirror the pipeline combs
    """: {
        coproc_response_cfg = coproc_response;
        if (coproc_force_disable || riscv_config.coproc_disable) {
            coproc_response_cfg = {*=0};
        }

        coproc_controls = {*=0};
        coproc_controls.dec_idecode_valid  = dec_state.valid;
        coproc_controls.dec_idecode        = dec_combs.idecode;
        coproc_controls.dec_to_alu_blocked = alu_combs.cannot_complete;
        coproc_controls.alu_rs1 = alu_combs.rs1;
        coproc_controls.alu_rs2 = alu_combs.rs2;
        coproc_controls.alu_flush_pipeline = alu_combs.flush_pipeline;
        coproc_controls.alu_cannot_start    = alu_combs.blocked_by_mem;
        coproc_controls.alu_cannot_complete = alu_combs.cannot_complete;
        if (coproc_force_disable || riscv_config.coproc_disable) {
            coproc_controls = {*=0};
        }
    }

    /*b Tracing */
    logging """
    """: {
        trace = {*=0};
        trace.instr_valid = alu_state.valid;
        trace.instr_pc    = alu_state.pc;
        trace.instruction = alu_state.debug_instruction;
        trace.rfw_retire     = rfw_state.valid;
        trace.rfw_data_valid = rfw_state.rd_written;
        trace.rfw_rd         = rfw_state.rd;
        trace.rfw_data       = rfw_state.mem_result;
        trace.branch_taken   = alu_combs.branch_taken || alu_combs.jalr;
        trace.trap           = alu_combs.trap;
        trace.branch_target  = alu_combs.next_pc;
    }

    /*b All done */
}

