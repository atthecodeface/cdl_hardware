/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   apb_target_led_ws2812.cdl
 * @brief  Simple APB target for driving a chain of Neopixels
 *
 * CDL implementation of a simple APB target to drive a chain of Neopixels.
 *
 */
/*a Includes
 */
include "apb.h"
include "leds.h"

/*a Types */
/*t t_apb_address
 *
 * APB address map, used to decode paddr
 */
typedef enum [5] {
    apb_address_config = 0   "Address of configuration register (number of LEDs and operating clock divisor)",
    apb_address_leds = 16    "Base address of 16 registers for RGB values of 16 LEDs", // 16 leds
} t_apb_address;

/*t t_access
 *
 * APB access that is in progress; a decode of psel and paddr
 */
typedef enum [3] {
    access_none           "No APB access",
    access_write_config   "APB write to the configuration register",
    access_read_config    "APB read of the configuration register",
    access_write_led      "APB write to an LED register, given by paddr[4;0]"
} t_access;

/*t t_rgb
 *
 * 24-bit RGB color
 *
 */
typedef struct
{
    bit[8] red    "Red component value";
    bit[8] green  "Green component value";
    bit[8] blue   "Blue component value";
} t_rgb;

/*t t_chain_state
 *
 * Clock divider and LED contents
 *
 */
typedef struct
{
    bit[8] divider_400ns  "Divider to generate approximately a 400ns period (e.g. for 50MHz, should be 400ns/20ns-1 = 19)";
    bit[4] last_led       "Last LED number, 0 (for 1 LED) to 15 (for 16 LEDs)";
} t_chain_state;

/*a Module */
module apb_target_led_ws2812( clock clk         "System clock",
                              input bit reset_n "Active low reset",

                              input  t_apb_request  apb_request  "APB request",
                              output t_apb_response apb_response "APB response",

                              input bit[8] divider_400ns_in "Default value for divider_400ns",

                              output bit led_chain
    )
"""
A simple module to drive a chain of Neopixel LEDs as an APB target.

The Neopixel LEDs are 24-bit RGB LEDs that are driven through a chain,
with a single control pin providing the information for the LEDs.

This module supports up to 16 LEDs in a chain, each with a 24-bit RGB
value. The chain must be configured with a clock divider (which is the
number of clock ticks required to generate a 400ns, approximately,
clock) and the number of LEDs in the chain.

The clock divider resets to 0, but whenever it is zero it resets to
the input value @a divider_400ns_in; hence it may be effectively
'hardwired'.

Once configured the LED colors can be individually written to
address-mapped registers. The LED chain automatically updates.

The configuration register is:

Bits     | Meaning
---------|---------
12;2     | zero
4;16     | last LED in the chain (0 for one LED, 15 for sixteen LEDs)
8;8      | zero
8;0      | clock divider to create a 400ns clock enable from system clock

Example divider values

System clock   |  Period | Divider
----------------------------------
50MHz          | 20ns    |   19
100MHz         | 10ns    |   39
20MHz          | 50ns    |   7


"""
{
    /*b Clock and reset */
    default clock clk;
    default reset active_low reset_n;

    /*b Decode APB interface */
    clocked t_access access=access_none   "Access being performed by APB";

    /*b LED chain state */
    clocked t_chain_state chain_state={*=0};
    clocked t_rgb[16] leds = {*=0};

    /*b LED chain signals */
    net  t_led_ws2812_request led_request;
    comb t_led_ws2812_data    led_data;
    net bit led_chain;

    /*b APB interface */
    apb_interface_logic """
    The APB interface is decoded to @a access when @p psel is asserted
    and @p penable is deasserted - this is the first cycle of an APB
    access. This permits the access type to be registered, so that the
    APB @p prdata can be driven from registers, and so that writes
    will occur correctly when @p penable is asserted.

    The APB read data @p prdata can then be generated based on @a
    access.
    """ : {
        /*b Decode access */
        access <= access_none;
        part_switch (bundle(apb_request.paddr[4],4b0)) {
        case apb_address_config: {
            access <= apb_request.pwrite ? access_write_config : access_read_config;
        }
        case apb_address_leds: {
            access <= apb_request.pwrite ? access_write_led : access_none;
        }
        }
        if (!apb_request.psel || apb_request.penable) {
            access <= access_none;
        }

        /*b Handle APB read data */
        apb_response = {*=0, pready=1};
        if (access==access_read_config) {
            apb_response.prdata = bundle( 12b0,
                                          chain_state.last_led,
                                          8b0,
                                          chain_state.divider_400ns
                );
        }

        /*b All done */
    }

    /*b Handle the led chain */
    led_chain_logic """
    The LED chain logic manages the configuration (last led and divider), the LED data values, and
    the LED chain.

    The divider is set to the input value if it is zeroed (as it would
    be at reset, or if configured with 0); the @a last_led must be
    configured.

    The LED data values are simply written.

    The LED chain uses the @a led_ws2812_chain module, which presents
    an LED number - in response the LED's color must be returned. This
    is done simply with a multiplexing of the LED values.

    """: {
        /*b Clock divider and last led - configuration */
        if (chain_state.divider_400ns==0) {
            chain_state.divider_400ns <= divider_400ns_in;
        }
        if (access==access_write_config) {
            chain_state.divider_400ns <= apb_request.pwdata[8; 0];
            chain_state.last_led      <= apb_request.pwdata[4;16];
        }

        /*b LED data values */
        if (access==access_write_led) {
            leds[apb_request.paddr[4;0]].red   <= apb_request.pwdata[8; 0];
            leds[apb_request.paddr[4;0]].green <= apb_request.pwdata[8; 8];
            leds[apb_request.paddr[4;0]].blue  <= apb_request.pwdata[8;16];
        }

        /*b LED chain */
        led_data = {*=0};
        if (led_request.ready) {
            led_data.red   = leds[led_request.led_number].red;
            led_data.green = leds[led_request.led_number].green;
            led_data.blue  = leds[led_request.led_number].blue;
            led_data.valid = 1;
            if (led_request.led_number[4;0] == chain_state.last_led) {
                led_data.last = 1;
            }
        }
        led_ws2812_chain leds( clk <- clk,
                               reset_n <= reset_n,
                               divider_400ns <= chain_state.divider_400ns,
                               led_request   => led_request,
                               led_data      <= led_data,
                               led_chain     => led_chain );
    }

    /*b Done
     */
}

/*a Editor preferences and notes
mode: c ***
c-basic-offset: 4 ***
c-default-style: (quote ((c-mode . "k&r") (c++-mode . "k&r"))) ***
outline-regexp: "/\\\*a\\\|[\t ]*\/\\\*[b-z][\t ]" ***
*/
