/** @copyright (C) 2019,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   tb_gbe.cdl
 * @brief  Testbench for gigabit ethernet with sgmii_gmii_gasket
 *
 */
/*a Includes */
include "types/ethernet.h"
include "networking/ethernet_modules.h"
include "networking/gmii_modules.h"

/*a External modules */
extern module axi4s32_master_slave( clock aclk,
                                    output t_axi4s32 master_axi4s,
                                    input bit      master_axi4s_tready,
                                    input t_tbi_valid tbi_tx "Optional TBI instead of SGMII",
                                    input bit[4] sgmii_txd,

                                    output t_tbi_valid tbi_rx "Optional TBI instead of SGMII",
                                    input t_axi4s32 slave_axi4s,
                                    output bit      slave_axi4s_tready,
                                    output t_timer_control rx_timer_control "Timer control for TX clock domain",
                                    output  t_sgmii_gasket_control sgmii_gasket_control "Control of gasket, on rx_clk",
                                    input t_sgmii_gasket_status  sgmii_gasket_status  "Status from gasket, on rx_clk",
                               
                                    output bit[32] sys_cfg
    )
{
    timing to   rising clock aclk master_axi4s_tready, tbi_tx, sgmii_txd;
    timing from rising clock aclk master_axi4s;
    timing from rising clock aclk slave_axi4s_tready, tbi_rx;
    timing to   rising clock aclk slave_axi4s;
    timing from rising clock aclk rx_timer_control;
    timing from rising clock aclk sys_cfg;
}

/*a Module */
module tb_gbe( clock clk,
                 input bit reset_n
)
{

    /*b Nets */
    net t_axi4s32 master_axi4s;
    net bit      master_axi4s_tready;

    net t_axi4s32 slave_axi4s;
    net bit      slave_axi4s_tready;
    net t_timer_control rx_timer_control;

    net t_gmii_tx gmii_tx;
    net bit gmii_tx_enable;

    net t_tbi_valid tbi_tx;
    net bit[4] sgmii_txd;
    net t_tbi_valid tbi_rx;
    net bit gmii_rx_enable;
    net t_gmii_rx gmii_rx;
    comb bit[4] sgmii_rxd;
    net bit[32] sys_cfg;
    net  t_sgmii_gasket_control sgmii_gasket_control "Control of gasket, on rx_clk";
    net t_sgmii_gasket_status   sgmii_gasket_status  "Status from gasket, on rx_clk";

    clocked clock clk reset active_low reset_n bit[16]         sgmii_stream=0;

    /*b Instantiations */
    instantiations: {
        axi4s32_master_slave th( aclk <- clk,
                                 master_axi4s => master_axi4s,
                                 master_axi4s_tready <= master_axi4s_tready,
                                 tbi_tx <= tbi_tx,
                                 sgmii_txd <= sgmii_txd,

                                 tbi_rx => tbi_rx,
                                 slave_axi4s <= slave_axi4s,
                                 slave_axi4s_tready => slave_axi4s_tready,
                                 rx_timer_control   => rx_timer_control,

                                 sgmii_gasket_control => sgmii_gasket_control,
                                 sgmii_gasket_status  <= sgmii_gasket_status,
                                 
                                 sys_cfg => sys_cfg );
        gbe_axi4s32 gbe( tx_aclk <- clk,
                     tx_areset_n <= reset_n,
                     tx_axi4s    <= master_axi4s,
                     tx_axi4s_tready => master_axi4s_tready,
                     gmii_tx_enable <= gmii_tx_enable,
                     gmii_tx        => gmii_tx,

                     rx_aclk <- clk,
                     rx_areset_n <= reset_n,
                     rx_axi4s => slave_axi4s,
                     rx_axi4s_tready <= slave_axi4s_tready,
                     gmii_rx_enable <= gmii_rx_enable,
                     gmii_rx <= gmii_rx,
                     rx_timer_control  <= rx_timer_control
            );
        sgmii_gmii_gasket sgg(tx_clk <- clk,
                              tx_clk_312_5 <- clk,
                              rx_clk <- clk,
                              rx_clk_312_5 <- clk,
                              tx_reset_n <= reset_n,
                              tx_reset_312_5_n <= reset_n,
                              rx_reset_n <= reset_n,
                              rx_reset_312_5_n <= reset_n,

                              gmii_tx <= gmii_tx,
                              gmii_tx_enable => gmii_tx_enable,
                              tbi_tx => tbi_tx,
                              sgmii_txd => sgmii_txd,

                              sgmii_rxd <= sgmii_rxd,
                              tbi_rx <= tbi_rx,
                              gmii_rx => gmii_rx,
                              gmii_rx_enable => gmii_rx_enable,

                              sgmii_gasket_control <= sgmii_gasket_control,
                              sgmii_gasket_status  => sgmii_gasket_status
            );
        sgmii_stream      <= sgmii_stream << 4;
        sgmii_stream[4;0] <= sgmii_txd;

        sgmii_rxd = sgmii_stream[4;1];
        if (sys_cfg[0]) {
            sgmii_rxd = sgmii_stream[4;0];
        }

        /*b All done */
    }

    /*b All done */
}

