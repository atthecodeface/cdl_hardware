/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   tb_riscv_i32_minimal.cdl
 * @brief  Testbench for minimal RISC-V
 *
 */

/*a Includes
 */
include "srams.h"
include "cpu/riscv/riscv.h"
include "cpu/riscv/riscv_modules.h"
include "types/apb.h"
include "apb/apb_targets.h"
include "apb/apb_masters.h"

/*a Constants
 */
constant integer i32c_force_disable=1;

/*a External modules */
extern module se_test_harness( clock clk, input bit a, output bit b )
{
    timing to rising clock clk a;
}

/*a Module
 */
module tb_riscv_i32_minimal( clock clk,
                             input bit reset_n
)
{

    /*b Nets
     */
    net t_sram_access_resp sram_access_resp;
    net t_sram_access_req sram_access_req;
    net t_riscv_mem_access_resp data_access_resp;
    net t_riscv_mem_access_req data_access_req;

    /*b State and comb
     */
    net bit[32] sram_ctrl;
    comb t_riscv_config riscv_config;
    default clock clk;
    default reset active_low reset_n;
    comb t_apb_request  th_apb_request;
    net t_apb_request   data_access_apb_request;
    net t_apb_request   mux_apb_request;
    comb t_apb_request  timer_apb_request;
    comb t_apb_request  sram_apb_request;
    net  t_apb_response timer_apb_response;
    net  t_apb_response sram_apb_response;
    comb t_apb_response mux_apb_response;
    net  t_apb_response data_access_apb_response;
    net  t_apb_response th_apb_response;
    comb t_timer_control timer_control;
    net t_timer_value timer_value;

    /*b Instantiate RISC-V
     */
    net t_riscv_i32_trace trace;
    comb t_riscv_irqs       irqs;
    riscv_instance: {
        riscv_config = {*=0};
        riscv_config.e32   = 0;
        riscv_config.i32c  = !i32c_force_disable;
        irqs = {*=0};
        irqs.mtip = timer_value.irq;
        th_apb_request = {*=0};
        riscv_i32_minimal_apb rv_apb( clk <- clk,
                                      reset_n <= reset_n,
                                      data_access_req  <= data_access_req,
                                      data_access_resp => data_access_resp,
                                      apb_request  => data_access_apb_request,
                                      apb_response <= data_access_apb_response );
    }
    apb_peripherals:
    {

        timer_control = {*=0};
        timer_control.enable_counter = 1;
        timer_control.fractional_adder = 2;
        timer_control.integer_adder    = 0;
        apb_master_mux apbmux( clk <- clk,
                               reset_n <= reset_n,
                               apb_request_0  <= data_access_apb_request,
                               apb_response_0 => data_access_apb_response,

                               apb_request_1 <= th_apb_request,
                               apb_response_1 => th_apb_response,

                               apb_request => mux_apb_request,
                               apb_response <= mux_apb_response
            );

        sram_apb_request  = mux_apb_request;
        timer_apb_request = mux_apb_request;

        timer_apb_request.psel = mux_apb_request.psel && (mux_apb_request.paddr[4;12]==0);
        sram_apb_request.psel  = mux_apb_request.psel && (mux_apb_request.paddr[4;12]==1);
        timer_apb_request.paddr = mux_apb_request.paddr >> 2;
        sram_apb_request.paddr = mux_apb_request.paddr >> 2;

        mux_apb_response = timer_apb_response;
        if (sram_apb_request.psel) { mux_apb_response = sram_apb_response; }

        apb_target_rv_timer timer( clk <- clk,
                                   reset_n <= reset_n,
                                   timer_control <= timer_control,
                                   apb_request  <= timer_apb_request,
                                   apb_response => timer_apb_response,
                                   timer_value => timer_value );

        apb_target_sram_interface sram_if( clk <- clk,
                                           reset_n <= reset_n,
                                           apb_request  <= sram_apb_request,
                                           apb_response => sram_apb_response,
                                           sram_ctrl    => sram_ctrl,
                                           sram_access_req => sram_access_req,
                                           sram_access_resp <= sram_access_resp );

        se_test_harness th( clk <- clk, a<=0 );
        
        riscv_i32_minimal dut( clk <- clk,
                               proc_reset_n <= reset_n & !sram_ctrl[0],
                               reset_n <= reset_n,
                               irqs <= irqs,
                               data_access_req => data_access_req,
                               data_access_resp <= data_access_resp,
                               sram_access_req <= sram_access_req,
                               sram_access_resp => sram_access_resp,
                               riscv_config <= riscv_config,
                               trace => trace
                         );
        riscv_i32_trace trace(clk <- clk,
                              reset_n <= reset_n,
                              trace <= trace );
    }
}
