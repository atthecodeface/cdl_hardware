/** Copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *   http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * @file  tb_csrs.cdl
 * @brief Testbench for CSR interfaces and bus
 *
 */
/*a Includes */
include "types/ps2.h"
include "input/ps2_modules.h"

/*a External modules */
extern module se_test_harness( clock clk,
                               input  t_ps2_pins ps2_in,
                               output t_ps2_pins ps2_out,
                               input t_ps2_rx_data ps2_rx_data,
                               input t_ps2_key_state ps2_key,
                               output bit[16] divider
    )
{
    timing from rising clock clk ps2_out;
    timing to   rising clock clk ps2_in;

    timing from rising clock clk divider;
    timing to   rising clock clk ps2_rx_data, ps2_key;
}

/*a Module */
module tb_input_devices( clock clk,
                         input bit reset_n
)
{

    /*b Nets */
    net t_ps2_pins ps2_in;
    net t_ps2_pins ps2_out;
    net t_ps2_rx_data ps2_rx_data;
    net bit[16] divider;
    net t_ps2_key_state  ps2_key;

    /*b Instantiations */
    instantiations: {
        se_test_harness th( clk <- clk,
                            ps2_in <= ps2_out,
                            ps2_out => ps2_in,
                            ps2_rx_data <= ps2_rx_data,
                            ps2_key <= ps2_key,
                            divider => divider );
        
        ps2_host ps2( clk <- clk,
                      reset_n <= reset_n,
                      ps2_in <= ps2_in,
                      ps2_out => ps2_out,
                      ps2_rx_data => ps2_rx_data,
                      divider <= divider );
        
        ps2_host_keyboard key_decode(clk <- clk,
                                     reset_n <= reset_n,
                                     ps2_rx_data <= ps2_rx_data,
                                     ps2_key     => ps2_key );
    }

    /*b All done */
}

/*a Editor preferences and notes
mode: c ***
c-basic-offset: 4 ***
c-default-style: (quote ((c-mode . "k&r") (c++-mode . "k&r"))) ***
outline-regexp: "/\\\*a\\\|[\t ]*\/\\\*[b-z][\t ]" ***
*/
