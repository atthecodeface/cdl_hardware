/** @copyright (C) 2018,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   apb_master_axi.cdl
 * @brief  AXI target to an APB master interface
 *
 * The AXI target supports 32-bit aligned 32-bit read/writes with full
 * byte enables only.
 * 
 * Other transactions return a slave error response
 *
 
 VGA CSRs are not being written to


 Add rotary inputs

 Add PS/2 inputs

 */

/*a Includes
 */
include "types/apb.h"
include "types/dprintf.h"
include "types/csr.h"
include "types/ps2.h"
include "types/led.h"
include "types/teletext.h"
include "types/video.h"
include "srams.h"
include "csr/csr_masters.h"
include "csr/csr_targets.h"
include "apb/apb_targets.h"
include "apb/apb_masters.h"
include "utils/dprintf_modules.h"
include "led/led_modules.h"
include "video/framebuffer_modules.h"
include "cpu/riscv/riscv_modules.h"
include "boards/de2.h"

/*a Constants */
constant integer num_dprintf_requesters=16;
constant bit[8] divider_400ns = 19; // 2.5MHz
constant bit[8] sr_divider    = 49; // 1MHz

/*a Modules */
/*m picorisc_de2
 *
 * Debug module for testing out HPS in the Cyclone-V FPGA
 *
 */
module picorisc_de2( clock clk,
                     input bit reset_n,

                     clock de2_audio_bclk,
                     input  t_de2_audio de2_audio_adc,
                     output t_de2_audio de2_audio_dac,

                     input  t_i2c de2_i2c_in,
                     output t_i2c de2_i2c_out,

                     input t_de2_inputs de2_inputs,
                     output t_de2_leds de2_leds,
                     output t_de2_lcd  de2_lcd,

                     input t_ps2_pins   de2_ps2_in,
                     output t_ps2_pins  de2_ps2_out,

                     clock de2_td_clk,
                     output bit de2_td_reset_n,
                     input t_adv7180 de2_td,

                     input t_uart_in   de2_uart_in,
                     output t_uart_out de2_uart_out,

                     clock de2_vga_clk,
                     input bit de2_vga_reset_n,
                     output t_adv7123 de2_vga,

                     clock de2_sdr_clk,
                     output t_sdram_16_12_2_out de2_sdr_out,
                     input  t_sdram_16_12_2_in  de2_sdr_in,

                     output t_asram_16_18_out de2_sram_out,
                     input  t_asram_16_18_in  de2_sram_in,

                     output t_flash_8_22_out de2_flash_out,
                     input  t_flash_8_22_in  de2_flash_in,

                     input t_de2_gpio de2_gpio_in
    )
{
    /*b Clock and reset */
    default clock clk;
    default reset active_low reset_n;
    /*b Nets */
    //net  t_apb_request riscv_apb_request;
    net  t_apb_request proc_apb_request;

    //net t_apb_request  rp_apb_request;
    comb t_apb_request  apb_request;
    comb bit[4]        apb_request_sel;
    comb t_apb_request timer_apb_request;
    comb t_apb_request dprintf_apb_request;
    comb t_apb_request csr_apb_request;
    comb t_apb_request rv_sram_apb_request;
    comb t_apb_request fb_sram_apb_request;
    comb t_apb_request ps2_apb_request;

    net t_apb_response  timer_apb_response;
    net t_apb_response  dprintf_apb_response;
    net t_apb_response  csr_apb_response;
    net t_apb_response  rv_sram_apb_response;
    net t_apb_response  fb_sram_apb_response;
    net t_apb_response  ps2_apb_response;
    comb t_apb_response apb_response;

    comb t_apb_response proc_apb_response;

    comb t_timer_control timer_control;
    net  t_timer_value timer_value;
    net bit[32] rv_sram_ctrl;
    net bit[32] fb_sram_ctrl;

    net  t_dprintf_req_4 apb_dprintf_req "Dprintf request from APB target";
    comb bit             apb_dprintf_ack "Ack for dprintf request from APB target";

    net bit[num_dprintf_requesters]                 dprintf_ack;
    clocked t_dprintf_req_4[num_dprintf_requesters] dprintf_req={*=0};
    net bit[num_dprintf_requesters-1]               mux_dprintf_ack "Ack for dprintf request after multiplexing";
    net t_dprintf_req_4[num_dprintf_requesters-1]   mux_dprintf_req "Dprintf request after multiplexing";
    net t_dprintf_byte dprintf_byte;

    net t_csr_request   csr_request;
    comb t_csr_response csr_response;
    clocked t_csr_response csr_response_r = {*=0};
    net t_csr_response tt_vga_framebuffer_csr_response;
    net t_csr_response timeout_csr_response;
    comb t_sram_access_req tt_display_sram_access_req;
    net t_video_bus vga_video_bus;

    clocked t_apb_processor_request  apb_processor_request={*=0};
    clocked bit apb_processor_completed = 0;
    net t_apb_processor_response  apb_processor_response;
    net t_apb_rom_request         apb_rom_request;
    net bit[40]                   apb_rom_data;

    /*
    comb t_riscv_config riscv_config;
    net t_riscv_i32_trace riscv_trace;
    comb t_riscv_irqs       irqs;
    net t_riscv_mem_access_req data_access_req;
    net t_riscv_mem_access_resp data_access_resp;
    */
    net t_sram_access_req  rv_sram_access_req;
    comb t_sram_access_resp rv_sram_access_resp;
    net t_sram_access_req  fb_sram_access_req;
    comb t_sram_access_resp fb_sram_access_resp;

    clocked bit[32] divider=0;
    clocked bit divider_reset=0;
    clocked bit[8]  seconds=0;
    clocked bit[32] counter=0;

    clocked t_ps2_pins       ps2_in = {*=-1};
    clocked t_ps2_pins  de2_ps2_out = {*=-1};
    net t_ps2_pins  ps2_out;

    net bit[7][6]de2_hex_leds;
//    clocked bit[32] riscv_last_pc=0;

    default clock de2_vga_clk;
    default reset active_low de2_vga_reset_n;
    clocked bit[4]  vga_vsync_counter=0;
    clocked bit[12] vga_hsync_counter=0;
    clocked t_adv7123 de2_vga={*=0};
    clocked bit[4] vga_seconds_sr = 0;
    clocked bit[32][4] vga_counters={*=0};

    /*b RISC-V */
    riscv_instance: {
        /*
        riscv_config = {*=0};
        riscv_config.e32   = 0;
        riscv_config.i32c  = 1;
        irqs = {*=0};
        irqs.mtip = timer_value.irq;

        riscv_i32_minimal riscv( clk <- clk,
                               proc_reset_n <= reset_n & rv_sram_ctrl[0],
                               reset_n <= reset_n,
                               irqs <= irqs,
                               data_access_req => data_access_req,
                               data_access_resp <= data_access_resp,
                               sram_access_req <= rv_sram_access_req,
                               sram_access_resp => rv_sram_access_resp,
                               riscv_config <= riscv_config,
                               trace => riscv_trace
                         );
        riscv_i32_trace trace(clk <- clk,
                              reset_n <= reset_n,
                              trace <= riscv_trace );

        riscv_i32_minimal_apb rv_apb( clk <- clk,
                                      reset_n <= reset_n,
                                      data_access_req  <= data_access_req,
                                      data_access_resp => data_access_resp,
                                      apb_request  => riscv_apb_request,
                                      apb_response <= riscv_apb_response );
    */
        timer_control = {*=0};
        timer_control.enable_counter = 1;
        timer_control.integer_adder = 20; // 50MHz
    }
    /*b APB processor */
    apb_master_instances: {
        apb_processor_request.address <= 0;
        apb_processor_request.valid   <= !apb_processor_completed;
        if (apb_processor_response.acknowledge) {
            apb_processor_request.valid   <= 0;
            apb_processor_completed <= 1;
        }

        apb_processor apbp( clk <- clk,
                            reset_n <= reset_n,

                            apb_processor_request <= apb_processor_request,
                            apb_processor_response => apb_processor_response,
                            apb_request   => proc_apb_request,
                            apb_response  <= proc_apb_response,
                            rom_request   => apb_rom_request,
                            rom_data      <= apb_rom_data );

        se_sram_srw_256x40 apb_rom(sram_clock <- clk,
                                   select <= apb_rom_request.enable,
                                   address <= apb_rom_request.address[8;0],
                                   read_not_write <= 1,
                                   write_data <= 0,
                                   data_out => apb_rom_data );

    }

    /*b APB master multiplexing and decode */
    apb_multiplexing_decode: {
        apb_request =  proc_apb_request;

        apb_request_sel = apb_request.paddr[4;16]; // 1MB of address space, top 4 bits as select
        timer_apb_request      = apb_request;
        dprintf_apb_request    = apb_request;
        csr_apb_request        = apb_request;
        rv_sram_apb_request    = apb_request;
        fb_sram_apb_request    = apb_request;
        ps2_apb_request        = apb_request;

        timer_apb_request.paddr      = apb_request.paddr >> 2;
        dprintf_apb_request.paddr    = apb_request.paddr >> 2;
        rv_sram_apb_request.paddr    = apb_request.paddr >> 2;
        fb_sram_apb_request.paddr    = apb_request.paddr >> 2;
        ps2_apb_request.paddr        = apb_request.paddr >> 2;

        timer_apb_request.psel       = apb_request.psel && (apb_request_sel==0);
        dprintf_apb_request.psel     = apb_request.psel && (apb_request_sel==2);
        csr_apb_request.psel         = apb_request.psel && (apb_request_sel==3);
        rv_sram_apb_request.psel     = apb_request.psel && (apb_request_sel==4);
        fb_sram_apb_request.psel     = apb_request.psel && (apb_request_sel==7);
        ps2_apb_request.psel         = apb_request.psel && (apb_request_sel==8);
        csr_apb_request.paddr[16;16] = bundle(12b0,apb_request.paddr[4;12]);
        csr_apb_request.paddr[16;0]  = bundle( 6b0,apb_request.paddr[10;2]);

        apb_response = timer_apb_response; // defaulting to timer is good - it is always ready even if not selected...
        if (apb_request_sel==2) { apb_response = dprintf_apb_response; }
        if (apb_request_sel==3) { apb_response = csr_apb_response; }
        if (apb_request_sel==4) { apb_response = rv_sram_apb_response; }
        if (apb_request_sel==7) { apb_response = fb_sram_apb_response; }
        if (apb_request_sel==8) { apb_response = ps2_apb_response; }
        proc_apb_response = apb_response;
    }

    /*b Dprintf requesting */
    dprintf_requesting : {
        for (i; num_dprintf_requesters) {
            if (dprintf_ack[i]) {
                dprintf_req[i].valid <= 0;
            }
        }
        dprintf_req[0] <= apb_dprintf_req;
        apb_dprintf_ack = dprintf_ack[0];

        if (apb_request.psel) {
            dprintf_req[6] <= {valid=1, address=240,
                    data_0=bundle(40h41_50_42_3a_80, 7b0,apb_request.pwrite, 16h_20_87), // APB:%x %08x %08x (pwrite paddr pwdata)
                    data_1=bundle(apb_request.paddr, 32h20000087),
                    data_2=bundle(apb_request.pwdata, 8hff, 24h0) };
        }
        if (csr_request.valid) {
            dprintf_req[7] <= {valid=1, address=280,
                    data_0=bundle(40h43_53_52_3a_80, 7b0,csr_request.read_not_write, 16h_20_83), // CSR:%x %04x %04x %08x (read_not_write select address data)
                    data_1=bundle(csr_request.select,  48h200000000083),
                    data_2=bundle(csr_request.address, 48h200000000087),
                    data_3=bundle(csr_request.data,    8hff, 24h0) };
        }
        if (rv_sram_access_req.valid) {
            dprintf_req[8] <= {valid=1, address=320,
                    data_0=bundle(40h53_52_4d_3a_83, 4b0,rv_sram_access_req.id,16h_20_80), // SRM:%x %x %08x %08x %x (id read_not_write address data be)
                    data_1=bundle(7b0,rv_sram_access_req.read_not_write,  56h20000000000087),
                    data_2=bundle(rv_sram_access_req.address,    32h20000087),
                    data_3=bundle(rv_sram_access_req.write_data[32;0], 16h2080, rv_sram_access_req.byte_enable, 8hff) };
        }
        if (divider_reset) {
            dprintf_req[11] <= {valid=1, address=440,
                    data_0=bundle(32h56_47_41_3a, 32h_00_00_00_87), // VGA:%08x %08x %08x (cnts0/1/2)
                    data_1=bundle(vga_counters[0], 32h20000087),
                    data_2=bundle(vga_counters[1], 32h20000087),
                    data_3=bundle(vga_counters[2], 8hff, 24h0) };
        }
    }

    /*b Dprintf multiplexing */
    dprintf_multiplexing """
    mux[n-2] = req[n-2] * req[n-1]
    mux[n-3] = req[n-2] * mux[n-2]
    mux[2]   = req[2] * mux[3]
    mux[1]   = req[1] * mux[2]
    mux[0]   = req[0] * mux[1]
    """: {
        dprintf_4_mux tdm_n( clk <- clk,
                             reset_n <= reset_n,
                             req_a <= dprintf_req[num_dprintf_requesters-2],
                             ack_a => dprintf_ack[num_dprintf_requesters-2],
                             req_b <= dprintf_req[num_dprintf_requesters-1],
                             ack_b => dprintf_ack[num_dprintf_requesters-1],
                             req => mux_dprintf_req[num_dprintf_requesters-2],
                             ack <= mux_dprintf_ack[num_dprintf_requesters-2] );

        for (i; num_dprintf_requesters-2) {
            dprintf_4_mux tdm[i]( clk <- clk, reset_n <= reset_n,
                                  req_a <= dprintf_req[i],
                                  ack_a => dprintf_ack[i],
                                  req_b <= mux_dprintf_req[i+1],
                                  ack_b => mux_dprintf_ack[i+1],
                                  req => mux_dprintf_req[i],
                                  ack <= mux_dprintf_ack[i] );
        }

    }

    /*b APB targets */
    apb_target_instances: {

        apb_target_sram_interface rv_sram_if( clk <- clk,
                                           reset_n <= reset_n,
                                           apb_request  <= rv_sram_apb_request,
                                           apb_response => rv_sram_apb_response,
                                           sram_ctrl    => rv_sram_ctrl,
                                           sram_access_req => rv_sram_access_req,
                                           sram_access_resp <= rv_sram_access_resp );

        apb_target_sram_interface fb_sram_if( clk <- clk,
                                           reset_n <= reset_n,
                                           apb_request  <= fb_sram_apb_request,
                                           apb_response => fb_sram_apb_response,
                                           sram_ctrl    => fb_sram_ctrl,
                                           sram_access_req => fb_sram_access_req,
                                           sram_access_resp <= fb_sram_access_resp );

        apb_target_dprintf apb_dprintf( clk <- clk,
                                    reset_n <= reset_n,
                                    apb_request  <= dprintf_apb_request,
                                    apb_response => dprintf_apb_response,
                                    dprintf_req => apb_dprintf_req,
                                    dprintf_ack <= apb_dprintf_ack );

        apb_target_rv_timer timer( clk <- clk,
                                   reset_n <= reset_n,
                                   timer_control <= timer_control,
                                   apb_request  <= timer_apb_request,
                                   apb_response => timer_apb_response,
                                   timer_value => timer_value );

        ps2_in <= de2_ps2_in;
        apb_target_ps2_host ps2_if( clk <- clk,
                                    reset_n <= reset_n,
                                    apb_request  <= ps2_apb_request,
                                    apb_response => ps2_apb_response,
                                    ps2_in  <= ps2_in,
                                    ps2_out => ps2_out );

        csr_master_apb master( clk <- clk,
                               reset_n <= reset_n,
                               apb_request <= csr_apb_request,
                               apb_response => csr_apb_response,
                               csr_request => csr_request,
                               csr_response <= csr_response_r );

    }

    /*b Dprintf/framebuffer */
    dprintf_framebuffer_instances: {
        dprintf dprintf( clk <- clk,
                         reset_n <= reset_n,
                         dprintf_req <= mux_dprintf_req[0],
                         dprintf_ack => mux_dprintf_ack[0],
                         dprintf_byte => dprintf_byte
            );

        tt_display_sram_access_req = {*=0,
                                      valid = dprintf_byte.valid,
                                      address = bundle(16b0, dprintf_byte.address),
                                      write_data = bundle(56b0, dprintf_byte.data) };

        fb_sram_access_resp = {*=0};
        fb_sram_access_resp.ack   = fb_sram_access_req.valid;
        fb_sram_access_resp.valid = fb_sram_access_req.valid;
        fb_sram_access_resp.id    = fb_sram_access_req.id;
        rv_sram_access_resp = {*=0};
        rv_sram_access_resp.ack   = rv_sram_access_req.valid;
        rv_sram_access_resp.valid = rv_sram_access_req.valid;
        rv_sram_access_resp.id    = rv_sram_access_req.id;

        framebuffer_teletext ftb_vga( csr_clk <- clk,
                                      sram_clk <- clk,
                                      video_clk <- de2_vga_clk,
                                      reset_n <= reset_n,
                                      video_bus => vga_video_bus,
                                      display_sram_write <= tt_display_sram_access_req,
                                      csr_select_in <= 16h4, // uses 2 selects
                                      csr_request <= csr_request,
                                      csr_response => tt_vga_framebuffer_csr_response
            );

        csr_target_timeout csr_timeout(clk <- clk,
                                       reset_n <= reset_n,
                                       csr_request <= csr_request,
                                       csr_response => timeout_csr_response,
                                       csr_timeout <= 16h100 );

        csr_response  = tt_vga_framebuffer_csr_response;
        csr_response |= timeout_csr_response;
        csr_response_r <= csr_response;

        de2_vga.hs <= 1;
        if (vga_hsync_counter!=0) {
            de2_vga.hs <= 0;
            vga_hsync_counter <= vga_hsync_counter-1;
        }
        if (vga_video_bus.hsync) {
            de2_vga.hs <= 0;
            vga_hsync_counter <= 110; // 128 for 64MHz officially, 96 for 25MHz
            de2_vga.vs <= 1;
            if (vga_vsync_counter!=0) {
                de2_vga.vs <= 0;
                vga_vsync_counter <= vga_vsync_counter-1;
            }
        }
        if (vga_video_bus.vsync) {
            de2_vga.vs <= 0;
            vga_vsync_counter <= 1;
        }
        
        de2_vga.blank_n <= vga_video_bus.display_enable;
        de2_vga.sync_n  <= de2_vga.vs & de2_vga.hs;
        if (de2_inputs.switches[9]) {
            de2_vga.sync_n  <= de2_inputs.switches[8];
        }
        de2_vga.red     <= bundle(vga_video_bus.red  [8;0],2b0);
        de2_vga.green   <= bundle(vga_video_bus.green[8;0],2b0);
        de2_vga.blue    <= bundle(vga_video_bus.blue [8;0],2b0);

        if (vga_video_bus.vsync) {
            vga_counters[0] <= vga_counters[0]+1;
        }
        if (vga_video_bus.hsync) {
            vga_counters[1] <= vga_counters[1]+1;
        }
        if (vga_video_bus.display_enable) {
            vga_counters[2] <= vga_counters[2]+1;
        }
        vga_seconds_sr <= bundle(seconds[0], vga_seconds_sr[3;1]);
        if (vga_seconds_sr[0]!=vga_seconds_sr[1]) {
            vga_counters[0] <= 0;
            vga_counters[1] <= 0;
            vga_counters[2] <= 0;
            vga_counters[3] <= 0;
        }

    }

    /*b Stub out unused outputs and all done */
    stubs : {
        divider <= divider+1;
        divider_reset <= 0;
        if (divider==50*1000*1000) {
            divider <= 0;
            divider_reset <= 1;
            seconds <= seconds + 1;
        }
        if (de2_inputs.switches[3;2]==0) {
            counter <= counter + 1;
        }
        if ((de2_inputs.switches[3;2]==1) && (mux_dprintf_req[0].valid)) {
            counter <= counter + 1;
        }
        if ((de2_inputs.switches[3;2]==2) && (mux_dprintf_ack[0])) {
            counter <= counter + 1;
        }
        if ((de2_inputs.switches[3;2]==3) && (apb_request.psel)) {
            counter <= counter + 1;
        }
        if ((de2_inputs.switches[3;2]==4) && (apb_processor_request.valid)) {
            counter <= counter + 1;
        }
        if ((de2_inputs.switches[3;2]==5) && (apb_processor_response.acknowledge)) {
            counter <= counter + 1;
        }
        if ((de2_inputs.switches[3;2]==6) && (tt_display_sram_access_req.valid)) {
            counter <= counter + 1;
        }

        for (i; 6) {
            led_seven_segment h[i](hex <= counter[4;4*i], leds=>de2_hex_leds[i] );
        }
        de2_leds = {*=0};
        de2_leds.ledr = counter[18;0];
        de2_leds.h0 = de2_hex_leds[0];
        de2_leds.h1 = de2_hex_leds[1];
        de2_leds.h2 = de2_hex_leds[2];
        de2_leds.h3 = de2_hex_leds[3];
        de2_leds.h4 = de2_hex_leds[4];
        de2_leds.h5 = de2_hex_leds[5];

        de2_ps2_out <= ps2_out;
    }
    /*b tieoffs */
    tieoffs: {
        de2_audio_dac = {*=0};
        de2_i2c_out = {*=1};
        de2_lcd = {*=0};
        de2_uart_out = {*=0};

        de2_td_reset_n = 0;
        de2_sdr_out = {*=0};
        de2_sram_out = {*=0};
        de2_flash_out = {*=0};
    }
}
