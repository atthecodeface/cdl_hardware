/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   riscv_i32_alu.cdl
 * @brief  ALU for i32 RISC-V implementation
 *
 * CDL implementation of RISC-V i32 ALU based on the RISC-V
 * specification v2.1.
 *
 */

/*a Includes
 */
include "cpu/riscv/riscv_pipeline_types.h"
include "cpu/riscv/riscv_internal_types.h"
include "cpu/riscv/riscv.h"

/*a Module
 */
module riscv_i32_pipeline_control_flow( input  t_riscv_pipeline_state     pipeline_state,
                                    input  t_riscv_pipeline_response  pipeline_response,
                                    output  t_riscv_pipeline_control  pipeline_control
    )
"""

"""
{
    code : {
        pipeline_control.valid = pipeline_state.valid;
        pipeline_control.fetch_action = pipeline_state.fetch_action;
        pipeline_control.fetch_pc = pipeline_state.fetch_pc;
        pipeline_control.mode = pipeline_state.mode;
        pipeline_control.error = pipeline_state.error;
        pipeline_control.tag = pipeline_state.tag;
        pipeline_control.halt = pipeline_state.halt;
        pipeline_control.interrupt_req = pipeline_state.interrupt_req;
        pipeline_control.interrupt_number = pipeline_state.interrupt_number;
        pipeline_control.ebreak_to_dbg = pipeline_state.ebreak_to_dbg;
        pipeline_control.interrupt_to_mode = pipeline_state.interrupt_to_mode;
        pipeline_control.instruction_data = pipeline_state.instruction_data;
        pipeline_control.instruction_debug = pipeline_state.instruction_debug;
        if (pipeline_response.rfw.valid) {
        pipeline_control.instruction_debug = pipeline_state.instruction_debug;
        }
    }
}
