/** Copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *   http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * @file   generic_valid_ack_mux.cdl
 * @brief  A generic valid/ack multiplexer to combine buses with valid/ack protocol
 *
 * CDL implementation of a module that takes a pair of input request
 * types, each of which has an individual @ack response signal, and it
 * combines them with a round-robin arbiter to a single request out.
 */
/*a Includes */

/*a Constants */

/*a Types */
/*t t_arbiter_state */
typedef struct {
    bit last_request_from_port_a "Asserted if the last request taken was from port A";
} t_arbiter_state;

/*t t_arbiter_combs */
typedef struct {
    bit new_request_permitted;
    bit take_req_a;
    bit take_req_b;
} t_arbiter_combs;

/*a Module
 */
module generic_valid_ack_mux( clock clk "Clock for data in and display SRAM write out",
                              input bit reset_n,
                              input gt_generic_valid_req req_a,
                              input gt_generic_valid_req req_b,
                              output bit ack_a,
                              output bit ack_b,
                              output gt_generic_valid_req req,
                              input bit ack
    )
"""
"""
{
    /*b State etc  */
    default reset active_low reset_n;
    default clock clk;

    clocked gt_generic_valid_req req={*=0};
    clocked bit ack_a=0;
    clocked bit ack_b=0;
    clocked t_arbiter_state arbiter_state={*=0};
    comb t_arbiter_combs arbiter_combs;

    /*b Arbiter logic */
    arbiter_logic """
    First determine if a new request may be presented.
    If it may, then chose one of the incoming requests, if either is valid.
    Else present NUL request.

    If a new request may not be presented then hold the output request
    stable and do not chose another request.
    """: {
        arbiter_combs.new_request_permitted = 0;
        if (!req.valid || ack) {
            arbiter_combs.new_request_permitted = 1;
        }

        arbiter_combs.take_req_a = 0;
        arbiter_combs.take_req_b = 0;
        if (arbiter_combs.new_request_permitted) {
            if ((req_a.valid && !ack_a) && (req_b.valid && !ack_b)) {
                arbiter_combs.take_req_a = !arbiter_state.last_request_from_port_a;
                arbiter_combs.take_req_b =  arbiter_state.last_request_from_port_a;
            } else {
                arbiter_combs.take_req_a = req_a.valid && !ack_a;
                arbiter_combs.take_req_b = req_b.valid && !ack_b;
            }
        }

        if (arbiter_combs.take_req_a) {
            arbiter_state.last_request_from_port_a <= 1;
        } elsif (arbiter_combs.take_req_b) {
            arbiter_state.last_request_from_port_a <= 0;
        }
    }
    
    /*b Input acknowledges and request output */
    input_ack_and_request_out_logic """
    Clear current request out if it is being acked.
    If taking a new request, then register that.
    Register the taking of a request as the ack to that requester.
    """: {
        ack_a <= arbiter_combs.take_req_a;
        ack_b <= arbiter_combs.take_req_b;

        if (ack) {
            req.valid <= 0;
        }
        if (arbiter_combs.take_req_a) {
            req <= req_a;
        }
        if (arbiter_combs.take_req_b) {
            req <= req_b;
        }

        /*b All done */
    }

    /*b All done */
}
