/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   tb_picoriscv.cdl
 * @brief  Testbench for Pico-RISC-V microcomputer
 *
 */

/*a Includes
 */
include "picoriscv.h"

/*a External modules */
extern module se_test_harness( clock clk,
                               input  t_apb_response apb_response,
                               output t_apb_request  apb_request
    )
{
    timing from rising clock clk apb_request;
    timing to   rising clock clk apb_response;
}


/*a Module
 */
module tb_picoriscv( clock clk,
                     input bit reset_n
)
{

    /*b Instantiate Pico-RISC-V microcomputer
     */
    net t_apb_request    th_apb_request;
    net t_apb_response   th_apb_response;
    net t_csr_request    csr_request;
    net t_csr_response   csr_response;
    comb t_prv_keyboard keyboard;
    riscv_instance: {
        keyboard = {*=0};
        se_test_harness th( clk <- clk,
                            apb_response <= th_apb_response,
                            apb_request  => th_apb_request );
        
        csr_master_apb master( clk <- clk,
                               reset_n <= reset_n,
                               apb_request <= th_apb_request,
                               apb_response => th_apb_response,
                               csr_request => csr_request,
                               csr_response <= csr_response );

        picoriscv dut(  clk <- clk,
                        reset_n <= reset_n,
                        video_clk <- clk,
                        video_reset_n <= reset_n,
                                         //video_bus,
                        keyboard <= keyboard,
                        csr_request <= csr_request,
                        csr_response => csr_response
                                    );
    }
}
