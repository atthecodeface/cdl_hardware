/** @copyright (C) 2019,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   apb_logging.cdl
 * @brief  Logging module for APB transactions
 *
 * This simple module provides a logging point for APB transactions, logging both
 * APB reads and writes separately.
 *
 * The module should be instantiated on an APB bus that the user wants
 * to have logged in CDL simulations
 *
 */
/*a Includes
 */
include "types/apb.h"

/*a Module
 */
module apb_logging( clock clk         "System clock",
                    input bit reset_n "Active low reset",

                    input t_apb_request  apb_request  "APB request",
                    input t_apb_response apb_response "APB response"
    )
"""
This simple module provides a logging point for APB transactions, logging both
APB reads and writes separately.

The module should be instantiated on an APB bus that the user wants
to have logged in CDL simulations
"""
{
    /*b Clock and reset */
    default clock clk;
    default reset active_low reset_n;

    /*b Logging */
    apb_logging """
    An APB transaction completes when @a psel, @a penable and @a pready are all high.
    Hence the @a pwdata and @prdata can be logged appropriately depending on @pwrite.
    """ : {
        /*b Logging */
        if (apb_request.psel && apb_request.penable && apb_response.pready) {
            if (apb_request.pwrite) {
                log("APB write",
                    "address", apb_request.paddr,
                    "data", apb_request.pwdata );
            } else {
                log("APB read",
                    "address", apb_request.paddr,
                    "data", apb_response.prdata );
            }
        }

        /*b All done */
    }

    /*b Done
     */
}
