/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   riscv_i32_trace.cdl
 * @brief  Instruction trace for RISC-V implementation
 *
 * CDL implementation of RISC-V instruction trace based on the RISC-V
 * specification v2.1.
 *
 */

/*a Includes
 */
include "cpu/riscv/riscv_internal_types.h"
include "cpu/riscv/riscv.h"

/*a Types
 */
typedef struct {
    bit[2]         must_be_ones "Bits that must be one for a valid RISCV I32 base instruction";
    bit            is_imm_op "Asserted if the instruction is an immediate operation";
    bit[5]         opc     "Opcode field from 32-bit instruction";
    bit[7]         funct7  "7-bit function field of instruction";
    bit[3]         funct3  "3-bit function field of instruction";
    t_riscv_word   imm_signed "Sign-extension word, basically instruction[31] replicated";
} t_combs;

/*a Module
 */
module riscv_i32_trace( clock clk            "Free-running clock",
                        input bit reset_n     "Active low reset",
                        input bit riscv_clk_enable "asserted if the RISC-V ticks on this edge",
                        input t_riscv_i32_trace trace "Trace signals"
)
"""
Trace instruction execution
"""
{

    default clock clk;
    default reset active_low reset_n;

    /*b Logging */
    logging """
    """ : {
        if (riscv_clk_enable) {
            if (trace.instr_valid) {
                log("PC",
                    "pc",trace.instr_pc,
                    "branch_taken",trace.branch_taken,
                    "branch_target",trace.branch_target,
                    "instr",trace.instruction.data);
                log("flow", "branch_taken", trace.branch_taken, "trap", trace.trap);
            }
            if (trace.rfw_retire) {
                log("retire", "rfw", trace.rfw_data_valid, "rd", trace.rfw_rd, "data", trace.rfw_data );
            }
        }
    }
    /*b All done */
}
