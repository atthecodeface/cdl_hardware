/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   tb_riscv_i32_minimal.cdl
 * @brief  Testbench for minimal RISC-V
 *
 */

/*a Includes
 */
include "srams.h"
include "riscv.h"
include "riscv_modules.h"
include "apb.h"
include "apb_peripherals.h"

/*a Constants
 */
constant integer i32c_force_disable=1;

/*a External modules */
extern module se_test_harness( clock clk, input bit a, output bit b )
{
    timing to rising clock clk a;
}

/*a Module
 */
module tb_riscv_i32_minimal( clock clk,
                             input bit reset_n
)
{

    /*b Nets
     */
    net t_sram_access_resp sram_access_resp;
    net t_riscv_mem_access_req data_access_req;

    /*b State and comb
     */
    comb t_sram_access_req sram_access_req;
    comb t_riscv_mem_access_resp data_access_resp;
    comb t_riscv_config riscv_config;
    default clock clk;
    default reset active_low reset_n;
    clocked t_apb_request apb_request={*=0};
    net t_apb_response apb_response;
    net bit[3] timer_equalled;

    /*b Instantiate RISC-V
     */
    net t_riscv_i32_trace trace;
    comb t_riscv_irqs       irqs;
    riscv_instance: {
        riscv_config = {*=0};
        riscv_config.e32   = 0;
        riscv_config.i32c  = !i32c_force_disable;
        irqs = {*=0};
        data_access_resp = {*=0};
        if (apb_request.psel) {
            data_access_resp.wait = 1;
            apb_request.penable <= 1;
            if (apb_request.penable && apb_response.pready) {
                apb_request.psel <= 0;
                apb_request.penable <= 0;
                data_access_resp.read_data = apb_response.prdata;
                data_access_resp.wait = 0;
            }
        } else {
            if (data_access_req.read_enable || data_access_req.write_enable) {
                data_access_resp.wait = 1;
                apb_request.psel <= 1;
                apb_request.penable <= 0;
                apb_request.paddr <= bundle(16b0,data_access_req.address[16;2]);
                apb_request.pwrite <= data_access_req.write_enable;
                apb_request.pwdata <= data_access_req.write_data;
            }
        }

        apb_target_timer timer( clk <- clk,
                                reset_n <= reset_n,
                                apb_request  <= apb_request,
                                apb_response => apb_response,
                                timer_equalled => timer_equalled );


        sram_access_req = {*=0};
        se_test_harness th( clk <- clk, a<=0 );
        
        riscv_i32_minimal dut( clk <- clk,
                               // add processor reset
                               reset_n <= reset_n,
                               irqs <= irqs,
                               data_access_req => data_access_req,
                               data_access_resp <= data_access_resp,
                               sram_access_req <= sram_access_req,
                               sram_access_resp => sram_access_resp,
                               riscv_config <= riscv_config,
                               trace => trace
                         );
        riscv_i32_trace trace(clk <- clk,
                              reset_n <= reset_n,
                              trace <= trace );
    }
}
