/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   tb_riscv_minimal.cdl
 * @brief  Testbench for minimal RISC-V
 *
 */

/*a Includes
 */
include "jtag.h"
include "apb.h"
include "apb_peripherals.h"

/*a External modules */
extern module se_test_harness( clock clk, output t_jtag jtag, input bit tdo )
{
    timing from rising clock clk jtag;
    timing to rising clock clk tdo;
}

/*a Module
 */
module tb_jtag_apb_timer( clock jtag_tck,
                          clock apb_clock,
                          input bit reset_n
)
{

    /*b Nets
     */
    net t_jtag jtag;
    net bit tdo;
    net bit[5]ir;
    net t_jtag_action dr_action;
    net bit[50]dr_in;
    net bit[50]dr_tdi_mask;
    net bit[50]dr_out;
    net t_apb_request apb_request;
    net t_apb_response apb_response;
    net bit[3] timer_equalled;

    /*b Instantiate APB timer
     */
    dut_instance: {
        se_test_harness th(clk <- jtag_tck, jtag=>jtag, tdo<=tdo);

        jtag_tap tap( jtag_tck <- jtag_tck,
                      reset_n <= reset_n,
                      jtag <= jtag,
                      tdo => tdo,

                      ir => ir,
                      dr_action => dr_action,
                      dr => dr_in,
                      dr_tdi_mask <= dr_tdi_mask,
                      dr_out <= dr_out );

        apb_target_timer timer( clk <- apb_clock,
                         reset_n <= reset_n,

                         apb_request <= apb_request,
                         apb_response => apb_response,

                         timer_equalled => timer_equalled
            );

        jtag_apb apb( jtag_tck <- jtag_tck,
                      reset_n <= reset_n,

                      ir <= ir,
                      dr_action <= dr_action,
                      dr_in <= dr_in,
                      dr_tdi_mask => dr_tdi_mask,
                      dr_out => dr_out,

                      apb_clock <- apb_clock,
                      apb_request => apb_request,
                      apb_response <= apb_response );
    }
}
