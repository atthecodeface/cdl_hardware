/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   apb_target_sram_interface.cdl
 * @brief  APB bus target to drive an SRAM read/write request
 *
 * CDL implementation of a simple APB target to interface to an SRAM
 * read/write request/response bus.
 *
 */
/*a Includes
 */
include "apb.h"
include "srams.h"

/*a Types */
/*t t_apb_address
 *
 * APB address map, used to decode paddr
 *
 * Each data or windowed access invokes a single sram access request
 *
 * This only supports 32-bit SRAM accesses.
 *
 */
typedef enum [8] {
    apb_address_address   = 0      "APB address for SRAM transaction request address",
    apb_address_data      = 1      "APB address for SRAM transaction request data; reading/writing makes an SRAM request occur",
    apb_address_control   = 2      "APB address for 32-bit SRAM control register",
    apb_address_data_inc  = 4      "Start of APB address range for data-with-autoincrement-of-address; reading/writing makes an SRAM request occur", // up to 128
    apb_address_windowed  = 128    "Start of APB address range for data addressed-by-window; reading/writing makes an SRAM request occur"
} t_apb_address;

/*t t_access
 *
 * APB access that is in progress; a decode of psel and paddr
 */
typedef enum [4] {
    access_none                   "No APB access",
    access_write_address          "Write SRAM address",
    access_read_address           "Read SRAM address",
    access_write_control          "Write SRAM control register",
    access_read_control           "Read SRAM control register",
    access_read_data              "Read SRAM data - by issuing SRAM transaction",
    access_read_data_inc          "Read SRAM data - by issuing SRAM transaction - and increment SRAM address",
    access_read_data_windowed     "Read SRAM data using paddr[7;0] as offset to address register - by issuing SRAM transaction",
    access_write_data             "Write SRAM data - by issuing SRAM transaction",
    access_write_data_inc         "Write SRAM data - by issuing SRAM transaction - and increment SRAM address",
    access_write_data_windowed    "Write SRAM data using paddr[7;0] as offset to address register - by issuing SRAM transaction",
} t_access;

/*t t_req_resp_state
 *
 * Timer comparator state; a 31-bit comparator with a single bit that
 * indicates if the timer value has incremented up to the comparator
 * value.
 */
typedef struct
{
    t_access access      "Access being performed";
    bit[32] address      "32 bit SRAM address";
    bit[32] control      "32 control bits to go to the SRAM";
    bit[32] data         "Data returned by SRAM read";
    bit     in_progress  "SRAM access in progress";
    bit     data_valid   "Asserted when SRAM read data is valid";
} t_req_resp_state;

/*a Module */
module apb_target_sram_interface( clock clk         "System clock",
                                  input bit reset_n "Active low reset",

                                  input  t_apb_request  apb_request  "APB request",
                                  output t_apb_response apb_response "APB response",

                                  output bit[32] sram_ctrl "SRAM control data, for whatever purpose",

                                  output t_sram_access_req  sram_access_req  "SRAM access request",
                                  input  t_sram_access_resp sram_access_resp "SRAM access response"
    )
"""
APB target peripheral that generates SRAM read/write requests

The module maintains a 32-bit SRAM address that is used in the
requests, which is a read/write register. There is also a 32-bit
control register, that can be used for any purpose by the client.

SRAM requests occur when the data register is accessed; it can be
accessed in one of three different ways. Firstly, it may be accessed
simply read/write, with either generating the appropriate SRAM request
to the address given by the SRAM address register. Secondly, it may be
accessed with a post-increment, where the SRAM address register value
is used as-is in the request, but it is incremented ready for a
subsequent transaction. Thirdly, it may be accessed 'windowed'; in
this manner the bottom 7 bits of the APB address are used in
conjunction with the top 25 bits of the SRAM address register to
generate the address for the SRAM request.

"""
{
    /*b Clock and reset */
    default clock clk;
    default reset active_low reset_n;

    /*b Decode APB interface */
    comb t_access access   "Access being performed by APB, combinatorial decode - only not none in first cycle";

    /*b Req/response state */
    clocked t_req_resp_state req_resp_state = {*=0};
    clocked t_sram_access_req  sram_access_req = {*=0, byte_enable=8h0f};

    /*b APB interface */
    apb_interface_logic """
    The APB interface is decoded to @a access when @p psel is asserted
    and @p penable is deasserted - this is the first cycle of an APB
    access. This permits the access type to be registered, so that the
    APB @p prdata can be driven from registers, and so that writes
    will occur correctly when @p penable is asserted.

    The APB read data @p prdata can then be generated based on @a
    access.
    """ : {
        /*b Decode access */
        access = access_none;
        if (apb_request.paddr[8;0] & apb_address_windowed) {
            access = apb_request.pwrite ? access_write_data_windowed : access_read_data_windowed;
        } else {
            part_switch (apb_request.paddr[7;0]) {
            case apb_address_address: {
                access = apb_request.pwrite ? access_write_address : access_read_address;
            }
            case apb_address_data: {
                access = apb_request.pwrite ? access_write_data : access_read_data;
            }
            case apb_address_control: {
                access = apb_request.pwrite ? access_write_control : access_read_control;
            }
            default: {
                access = apb_request.pwrite ? access_write_data_inc : access_read_data_inc;
            }
            }
        }
        if (!apb_request.psel || apb_request.penable) {
            access = access_none;
        }

        /*b Handle APB read data */
        sram_ctrl = req_resp_state.control;
        apb_response = {*=0, pready=1};
        part_switch (req_resp_state.access) {
        case access_read_address: {
            apb_response.prdata = req_resp_state.address;
        }
        case access_read_control: {
            apb_response.prdata = req_resp_state.control;
        }
        case access_read_data, access_read_data_inc, access_read_data_windowed: {
            apb_response.prdata = req_resp_state.data;
            apb_response.pready = req_resp_state.data_valid;
        }
        case access_write_data, access_write_data_inc, access_write_data_windowed: {
            apb_response.pready = !req_resp_state.in_progress;
        }
        }

        /*b All done */
    }

    /*b Handle SRAM requests */
    sram_request_logic """
    While an SRAM request is in progress the APB side is ignored; it
    should be held as busy. Hence an acknowledged valid request can be
    removed, and a valid SRAM response completes the SRAM request in
    progress.

    If an SRAM request is not in progress then one may be started,
    depending on the APB access being presented.
    """: {
        sram_access_req.id <= 0;
        sram_access_req.byte_enable <= 8h0f;
        if (req_resp_state.in_progress) {
            if (sram_access_req.valid && sram_access_resp.ack) {
                sram_access_req.valid <= 0;
            }
            if (sram_access_resp.valid) {
                req_resp_state.in_progress <= 0;
                req_resp_state.data <= sram_access_resp.data[32;0];
                req_resp_state.data_valid <= 1;
            }
        } else {
            if (access!=access_none) {
                req_resp_state.access <= access;
            }
            part_switch (access) {
            case access_write_address: {
                req_resp_state.address <= apb_request.pwdata;
            }
            case access_write_control: {
                req_resp_state.control <= apb_request.pwdata;
            }
            case access_read_data, access_read_data_inc, access_read_data_windowed: {
                sram_access_req.valid <= 1;
                sram_access_req.read_not_write <= 1;
                sram_access_req.address <= req_resp_state.address;
                req_resp_state.in_progress <= 1;
                req_resp_state.data_valid <= 0;
            }
            case access_write_data, access_write_data_inc, access_write_data_windowed: {
                sram_access_req.valid <= 1;
                sram_access_req.read_not_write <= 0;
                sram_access_req.address <= req_resp_state.address;
                sram_access_req.write_data <= bundle(32b0, apb_request.pwdata);
                req_resp_state.in_progress <= 1;
                req_resp_state.data_valid <= 0;
            }
            }
            if ( (access == access_write_data_windowed) || (access == access_read_data_windowed)) {
                sram_access_req.address[7;0] <= apb_request.paddr[7;0];
            }
            if ( (access == access_write_data_inc) || (access == access_read_data_inc)) {
                req_resp_state.address <= req_resp_state.address + 1;
            }
        }


    }

    /*b Done
     */
}

/*a Editor preferences and notes
mode: c ***
c-basic-offset: 4 ***
c-default-style: (quote ((c-mode . "k&r") (c++-mode . "k&r"))) ***
outline-regexp: "/\\\*a\\\|[\t ]*\/\\\*[b-z][\t ]" ***
*/
