/** @copyright (C) 2016-2017,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   riscv_minimal.cdl
 * @brief  Minimal RISC-V implementation ported to CDL
 *
 * CDL implementation of minimal RISC-V teaching implementation
 *
 * This is a two-stage pipeline implementation, with instruction fetch
 * of the next PC occuring simultaneously with the decode, register
 * read, ALU, data read/write request, data read memory access, and
 * register update.
 *
 * The instruction memory request, then, becomes valid dependent on
 * the decode of the registered instruction last fetched. For most
 * branches this requires only a small amount of logic, but for
 * jump-and-link-register instructions (which uses the full ALU
 * result) this may take a considerable amount of gates to determine
 * the correct branch target and hence next instruction fetch.  Hence
 * the instruction memory request is valid after a considerable delay
 * from the start of the cycle.
 *
 * The return value from the instruction memory request must be valid
 * before the end of the cycle.
 *
 * Any instruction memory implementation must start its access well
 * after the CPU clock edge, , as the request is valid after the CPU
 * clock edge; the resultant read data delay (from the clock edge)
 * then has to be factored in to determine when the next CPU clock
 * edge can occur. Hence it may be sensible to use a double speed
 * clock (e.g. 'fast_clk') to generate CPU clock edges (every other
 * fast_clk edge) and SRAM access clock edges (for a synchronous
 * memory) on the intervening fast_clk edges.
 *
 * The data memory request becomes valid, again, a fair time after the
 * CPU clock edge, as it requires instruction decode, register fetch,
 * and ALU operation to occur prior to the memory address being valid.
 *
 * The data memory response must be valid (for read data!) in the same
 * CPU cycle, as the returning data has to be rotated to the correct
 * byte lanes and prepared for the register file write.
 *
 * Hence a data memory implementation can be similar to that proposed
 * for the instruction memory - that is, accesses start on a memory
 * clock edge that is in the middle of a CPU clock edge, by using a
 * fast_clk.
 *
 */

/*a Includes
 */
include "cpu/riscv/riscv_internal_types.h"

/*a Types
 */
/*t t_ifetch_combs
 *
 * Combinatorials for the instruction fetch
 */
typedef struct {
    bit[32] pc_plus_4;
    bit[32] pc_plus_2;
    bit[32] pc_plus_inst;
} t_ifetch_combs;

/*a Module
 */
module riscv_i32_pipeline_control_fetch_req( input t_riscv_pipeline_control    pipeline_control,
                                             input t_riscv_pipeline_response   pipeline_response,
                                             output t_riscv_fetch_req          ifetch_req
)
{
    comb t_ifetch_combs ifetch_combs;
    /*b Pipeline control
     */
    pipeline_control_logic
    """
    The instruction fetch request derives from the
    decode/execute stage (the instruction address that is required
    next) and presents that to the outside world.

    This request may be for any 16-bit aligned address, and two
    successive 16-bit words from that request must be presented,
    aligned to bit 0.

    If the decode/execute stage is invalid (i.e. it does not have a
    valid instruction to decode) then the current PC is requested.
    """:
    {
        ifetch_req                 = {*=0};
        ifetch_req.valid           = 0;
        ifetch_req.sequential      = 0;
        ifetch_req.address         = pipeline_control.start_pc;
        ifetch_combs.pc_plus_4     = pipeline_response.decode.pc + 4;
        ifetch_combs.pc_plus_2     = pipeline_response.decode.pc + 2;
        ifetch_combs.pc_plus_inst  = ifetch_combs.pc_plus_4;
        if (pipeline_response.decode.is_compressed) {
            ifetch_combs.pc_plus_inst = ifetch_combs.pc_plus_2;
        }

        if (pipeline_control.fetch_action == rv_pc_fetch_action_restart_at_pc) {
            ifetch_req.valid   = 1;
            ifetch_req.address         = pipeline_control.start_pc;
        } elsif (pipeline_control.fetch_action == rv_pc_fetch_action_continue_fetching) {
            ifetch_req.valid = 1;
            ifetch_req.sequential = 1;
            if (pipeline_response.exec.action == rv_pipe_epc_flush) {
                ifetch_req.address = pipeline_response.exec.flush_target;
                ifetch_req.sequential = 0;
            } elsif (pipeline_response.decode.action==rv_pipe_dpc_flush) { // cannot happen on one-stage pipeline
            } elsif (pipeline_response.decode.action==rv_pipe_dpc_ret)   { // cannot happen on one-stage pipeline
            } elsif (pipeline_response.decode.action==rv_pipe_dpc_predict_branch) {  // cannot happen on one-stage pipeline
            } elsif (pipeline_response.decode.action==rv_pipe_dpc_sequential) {
                ifetch_req.sequential = 1;
                ifetch_req.address = ifetch_combs.pc_plus_inst;
            }
            if (pipeline_response.exec.trap.valid) { // vector interrupts if required
                ifetch_req.address = bundle(pipeline_response.exec.mtvec.base, 2b0);
                ifetch_req.sequential = 0;
                // flush if pipeline exists
            }
        }
    }
}
