/** @copyright (C) 2018,  Gavin J Stark.  All rights reserved.
 *
 * @copyright
 *    Licensed under the Apache License, Version 2.0 (the "License");
 *    you may not use this file except in compliance with the License.
 *    You may obtain a copy of the License at
 *     http://www.apache.org/licenses/LICENSE-2.0.
 *   Unless required by applicable law or agreed to in writing, software
 *   distributed under the License is distributed on an "AS IS" BASIS,
 *   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 *   See the License for the specific language governing permissions and
 *   limitations under the License.
 *
 * @file   riscv_i32_fetch_debug.cdl
 * @brief  Instruction fetch interposer for debug
 *
 * CDL implementation of RISC-V i32 instruction fetch interposer designed
 * to work with the pipeline and associated stateful debug modules
 *
 */

/*a Includes
 */
include "cpu/riscv/riscv_internal_types.h"
include "cpu/riscv/riscv.h"

/*a Types
 */
/*a Module
 */
module riscv_i32_fetch_debug( input  t_riscv_fetch_req  pipeline_ifetch_req,
                              output t_riscv_fetch_resp pipeline_ifetch_resp,
                              input  t_riscv_i32_trace pipeline_trace,
                              input  t_riscv_pipeline_debug_control debug_control,
                              output t_riscv_pipeline_debug_control debug_response,
                              output t_riscv_fetch_req  ifetch_req,
                              input  t_riscv_fetch_resp ifetch_resp
    )
"""

"""
{

    /*b Signals - just the combs */
    //comb t_fetch_debug_combs fetch_debug_combs      "Combinatorials used in the module, not exported as the decode";

    /*b FETCH_DEBUG operation */
    fetch_debug_operation """
    """ : {
        ifetch_req = pipeline_ifetch_req;
        pipeline_ifetch_resp = ifetch_resp;

        debug_response = {*=0};

        /*b All done */
    }

    /*b All done */
}
